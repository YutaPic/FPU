`default_nettype none
`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Yuta Fukushima
// 
// Create Date: 2020/10/31
// Design Name: fsqrt_table
// Module Name: fsqrt_const_table, fsqrt_grad_table
// Project Name: C&P
// Target Devices: KCU105
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
//////////////////////////////////////////////////////////////////////////////////
module fsqrt_const_table (
    input wire clk, 
    input wire [9:0] addr,
    output reg [22:0] con);

    reg [22:0] RAM [1023:0];
    always @(posedge clk)
        con <= RAM[addr];
    initial begin
        RAM[0] = 23'h3504f4;
        RAM[1] = 23'h35322f;
        RAM[2] = 23'h355f60;
        RAM[3] = 23'h358c85;
        RAM[4] = 23'h35b99f;
        RAM[5] = 23'h35e6ae;
        RAM[6] = 23'h3613b1;
        RAM[7] = 23'h3640a9;
        RAM[8] = 23'h366d96;
        RAM[9] = 23'h369a79;
        RAM[10] = 23'h36c750;
        RAM[11] = 23'h36f41c;
        RAM[12] = 23'h3720de;
        RAM[13] = 23'h374d94;
        RAM[14] = 23'h377a3f;
        RAM[15] = 23'h37a6e0;
        RAM[16] = 23'h37d376;
        RAM[17] = 23'h380001;
        RAM[18] = 23'h382c81;
        RAM[19] = 23'h3858f6;
        RAM[20] = 23'h388561;
        RAM[21] = 23'h38b1c1;
        RAM[22] = 23'h38de17;
        RAM[23] = 23'h390a61;
        RAM[24] = 23'h3936a2;
        RAM[25] = 23'h3962d7;
        RAM[26] = 23'h398f02;
        RAM[27] = 23'h39bb22;
        RAM[28] = 23'h39e739;
        RAM[29] = 23'h3a1345;
        RAM[30] = 23'h3a3f46;
        RAM[31] = 23'h3a6b3d;
        RAM[32] = 23'h3a9729;
        RAM[33] = 23'h3ac30b;
        RAM[34] = 23'h3aeee3;
        RAM[35] = 23'h3b1ab1;
        RAM[36] = 23'h3b4674;
        RAM[37] = 23'h3b722d;
        RAM[38] = 23'h3b9ddc;
        RAM[39] = 23'h3bc981;
        RAM[40] = 23'h3bf51b;
        RAM[41] = 23'h3c20ac;
        RAM[42] = 23'h3c4c33;
        RAM[43] = 23'h3c77af;
        RAM[44] = 23'h3ca321;
        RAM[45] = 23'h3cce8a;
        RAM[46] = 23'h3cf9e8;
        RAM[47] = 23'h3d253d;
        RAM[48] = 23'h3d5087;
        RAM[49] = 23'h3d7bc8;
        RAM[50] = 23'h3da6ff;
        RAM[51] = 23'h3dd22c;
        RAM[52] = 23'h3dfd4f;
        RAM[53] = 23'h3e2868;
        RAM[54] = 23'h3e5378;
        RAM[55] = 23'h3e7e7d;
        RAM[56] = 23'h3ea97a;
        RAM[57] = 23'h3ed46c;
        RAM[58] = 23'h3eff55;
        RAM[59] = 23'h3f2a34;
        RAM[60] = 23'h3f5509;
        RAM[61] = 23'h3f7fd6;
        RAM[62] = 23'h3faa98;
        RAM[63] = 23'h3fd551;
        RAM[64] = 23'h400000;
        RAM[65] = 23'h402aa7;
        RAM[66] = 23'h405543;
        RAM[67] = 23'h407fd6;
        RAM[68] = 23'h40aa5f;
        RAM[69] = 23'h40d4e0;
        RAM[70] = 23'h40ff56;
        RAM[71] = 23'h4129c4;
        RAM[72] = 23'h415429;
        RAM[73] = 23'h417e84;
        RAM[74] = 23'h41a8d5;
        RAM[75] = 23'h41d31e;
        RAM[76] = 23'h41fd5d;
        RAM[77] = 23'h422793;
        RAM[78] = 23'h4251bf;
        RAM[79] = 23'h427be4;
        RAM[80] = 23'h42a5fe;
        RAM[81] = 23'h42d010;
        RAM[82] = 23'h42fa18;
        RAM[83] = 23'h432418;
        RAM[84] = 23'h434e0e;
        RAM[85] = 23'h4377fb;
        RAM[86] = 23'h43a1e0;
        RAM[87] = 23'h43cbbb;
        RAM[88] = 23'h43f58d;
        RAM[89] = 23'h441f57;
        RAM[90] = 23'h444917;
        RAM[91] = 23'h4472cf;
        RAM[92] = 23'h449c7e;
        RAM[93] = 23'h44c624;
        RAM[94] = 23'h44efc1;
        RAM[95] = 23'h451956;
        RAM[96] = 23'h4542e2;
        RAM[97] = 23'h456c64;
        RAM[98] = 23'h4595de;
        RAM[99] = 23'h45bf51;
        RAM[100] = 23'h45e8b9;
        RAM[101] = 23'h461219;
        RAM[102] = 23'h463b71;
        RAM[103] = 23'h4664c0;
        RAM[104] = 23'h468e06;
        RAM[105] = 23'h46b744;
        RAM[106] = 23'h46e07a;
        RAM[107] = 23'h4709a6;
        RAM[108] = 23'h4732ca;
        RAM[109] = 23'h475be6;
        RAM[110] = 23'h4784f9;
        RAM[111] = 23'h47ae04;
        RAM[112] = 23'h47d706;
        RAM[113] = 23'h480000;
        RAM[114] = 23'h4828f2;
        RAM[115] = 23'h4851db;
        RAM[116] = 23'h487abc;
        RAM[117] = 23'h48a395;
        RAM[118] = 23'h48cc65;
        RAM[119] = 23'h48f52d;
        RAM[120] = 23'h491dec;
        RAM[121] = 23'h4946a3;
        RAM[122] = 23'h496f53;
        RAM[123] = 23'h4997fa;
        RAM[124] = 23'h49c099;
        RAM[125] = 23'h49e92f;
        RAM[126] = 23'h4a11be;
        RAM[127] = 23'h4a3a44;
        RAM[128] = 23'h4a62c2;
        RAM[129] = 23'h4a8b38;
        RAM[130] = 23'h4ab3a6;
        RAM[131] = 23'h4adc0c;
        RAM[132] = 23'h4b046a;
        RAM[133] = 23'h4b2cc0;
        RAM[134] = 23'h4b550e;
        RAM[135] = 23'h4b7d54;
        RAM[136] = 23'h4ba592;
        RAM[137] = 23'h4bcdc8;
        RAM[138] = 23'h4bf5f6;
        RAM[139] = 23'h4c1e1c;
        RAM[140] = 23'h4c463b;
        RAM[141] = 23'h4c6e51;
        RAM[142] = 23'h4c9660;
        RAM[143] = 23'h4cbe66;
        RAM[144] = 23'h4ce665;
        RAM[145] = 23'h4d0e5c;
        RAM[146] = 23'h4d364b;
        RAM[147] = 23'h4d5e33;
        RAM[148] = 23'h4d8613;
        RAM[149] = 23'h4dadeb;
        RAM[150] = 23'h4dd5bc;
        RAM[151] = 23'h4dfd84;
        RAM[152] = 23'h4e2545;
        RAM[153] = 23'h4e4cfe;
        RAM[154] = 23'h4e74b0;
        RAM[155] = 23'h4e9c5a;
        RAM[156] = 23'h4ec3fd;
        RAM[157] = 23'h4eeb98;
        RAM[158] = 23'h4f132b;
        RAM[159] = 23'h4f3ab7;
        RAM[160] = 23'h4f623b;
        RAM[161] = 23'h4f89b7;
        RAM[162] = 23'h4fb12c;
        RAM[163] = 23'h4fd89a;
        RAM[164] = 23'h500000;
        RAM[165] = 23'h50275f;
        RAM[166] = 23'h504eb6;
        RAM[167] = 23'h507606;
        RAM[168] = 23'h509d4f;
        RAM[169] = 23'h50c490;
        RAM[170] = 23'h50ebca;
        RAM[171] = 23'h5112fc;
        RAM[172] = 23'h513a27;
        RAM[173] = 23'h51614b;
        RAM[174] = 23'h518866;
        RAM[175] = 23'h51af7c;
        RAM[176] = 23'h51d68a;
        RAM[177] = 23'h51fd90;
        RAM[178] = 23'h52248f;
        RAM[179] = 23'h524b88;
        RAM[180] = 23'h527278;
        RAM[181] = 23'h529961;
        RAM[182] = 23'h52c044;
        RAM[183] = 23'h52e71f;
        RAM[184] = 23'h530df4;
        RAM[185] = 23'h5334c0;
        RAM[186] = 23'h535b87;
        RAM[187] = 23'h538245;
        RAM[188] = 23'h53a8fd;
        RAM[189] = 23'h53cfae;
        RAM[190] = 23'h53f657;
        RAM[191] = 23'h541cf9;
        RAM[192] = 23'h544395;
        RAM[193] = 23'h546a29;
        RAM[194] = 23'h5490b7;
        RAM[195] = 23'h54b73d;
        RAM[196] = 23'h54ddbd;
        RAM[197] = 23'h550435;
        RAM[198] = 23'h552aa7;
        RAM[199] = 23'h555111;
        RAM[200] = 23'h557775;
        RAM[201] = 23'h559dd2;
        RAM[202] = 23'h55c427;
        RAM[203] = 23'h55ea76;
        RAM[204] = 23'h5610bf;
        RAM[205] = 23'h563700;
        RAM[206] = 23'h565d3b;
        RAM[207] = 23'h56836f;
        RAM[208] = 23'h56a99c;
        RAM[209] = 23'h56cfc1;
        RAM[210] = 23'h56f5e1;
        RAM[211] = 23'h571bfa;
        RAM[212] = 23'h57420c;
        RAM[213] = 23'h576817;
        RAM[214] = 23'h578e1b;
        RAM[215] = 23'h57b419;
        RAM[216] = 23'h57da10;
        RAM[217] = 23'h580000;
        RAM[218] = 23'h5825ea;
        RAM[219] = 23'h584bcd;
        RAM[220] = 23'h5871aa;
        RAM[221] = 23'h58977f;
        RAM[222] = 23'h58bd4f;
        RAM[223] = 23'h58e317;
        RAM[224] = 23'h5908d9;
        RAM[225] = 23'h592e95;
        RAM[226] = 23'h59544a;
        RAM[227] = 23'h5979f8;
        RAM[228] = 23'h599fa0;
        RAM[229] = 23'h59c541;
        RAM[230] = 23'h59eadc;
        RAM[231] = 23'h5a1070;
        RAM[232] = 23'h5a35fe;
        RAM[233] = 23'h5a5b86;
        RAM[234] = 23'h5a8107;
        RAM[235] = 23'h5aa681;
        RAM[236] = 23'h5acbf5;
        RAM[237] = 23'h5af163;
        RAM[238] = 23'h5b16cb;
        RAM[239] = 23'h5b3c2b;
        RAM[240] = 23'h5b6186;
        RAM[241] = 23'h5b86da;
        RAM[242] = 23'h5bac28;
        RAM[243] = 23'h5bd170;
        RAM[244] = 23'h5bf6b1;
        RAM[245] = 23'h5c1bec;
        RAM[246] = 23'h5c4121;
        RAM[247] = 23'h5c664e;
        RAM[248] = 23'h5c8b77;
        RAM[249] = 23'h5cb099;
        RAM[250] = 23'h5cd5b4;
        RAM[251] = 23'h5cfac9;
        RAM[252] = 23'h5d1fd9;
        RAM[253] = 23'h5d44e1;
        RAM[254] = 23'h5d69e5;
        RAM[255] = 23'h5d8ee1;
        RAM[256] = 23'h5db3d7;
        RAM[257] = 23'h5dd8c8;
        RAM[258] = 23'h5dfdb2;
        RAM[259] = 23'h5e2296;
        RAM[260] = 23'h5e4773;
        RAM[261] = 23'h5e6c4b;
        RAM[262] = 23'h5e911d;
        RAM[263] = 23'h5eb5e8;
        RAM[264] = 23'h5edaae;
        RAM[265] = 23'h5eff6d;
        RAM[266] = 23'h5f2427;
        RAM[267] = 23'h5f48da;
        RAM[268] = 23'h5f6d87;
        RAM[269] = 23'h5f922e;
        RAM[270] = 23'h5fb6cf;
        RAM[271] = 23'h5fdb6b;
        RAM[272] = 23'h600000;
        RAM[273] = 23'h602490;
        RAM[274] = 23'h604919;
        RAM[275] = 23'h606d9c;
        RAM[276] = 23'h609219;
        RAM[277] = 23'h60b691;
        RAM[278] = 23'h60db03;
        RAM[279] = 23'h60ff6e;
        RAM[280] = 23'h6123d4;
        RAM[281] = 23'h614834;
        RAM[282] = 23'h616c8e;
        RAM[283] = 23'h6190e3;
        RAM[284] = 23'h61b531;
        RAM[285] = 23'h61d97a;
        RAM[286] = 23'h61fdbc;
        RAM[287] = 23'h6221f9;
        RAM[288] = 23'h624630;
        RAM[289] = 23'h626a61;
        RAM[290] = 23'h628e8d;
        RAM[291] = 23'h62b2b2;
        RAM[292] = 23'h62d6d3;
        RAM[293] = 23'h62faec;
        RAM[294] = 23'h631f01;
        RAM[295] = 23'h634310;
        RAM[296] = 23'h636719;
        RAM[297] = 23'h638b1c;
        RAM[298] = 23'h63af1a;
        RAM[299] = 23'h63d312;
        RAM[300] = 23'h63f705;
        RAM[301] = 23'h641af1;
        RAM[302] = 23'h643ed8;
        RAM[303] = 23'h6462b9;
        RAM[304] = 23'h648695;
        RAM[305] = 23'h64aa6b;
        RAM[306] = 23'h64ce3c;
        RAM[307] = 23'h64f206;
        RAM[308] = 23'h6515cc;
        RAM[309] = 23'h65398b;
        RAM[310] = 23'h655d46;
        RAM[311] = 23'h6580fa;
        RAM[312] = 23'h65a4a9;
        RAM[313] = 23'h65c852;
        RAM[314] = 23'h65ebf6;
        RAM[315] = 23'h660f95;
        RAM[316] = 23'h66332e;
        RAM[317] = 23'h6656c1;
        RAM[318] = 23'h667a4e;
        RAM[319] = 23'h669dd7;
        RAM[320] = 23'h66c15a;
        RAM[321] = 23'h66e4d8;
        RAM[322] = 23'h67084f;
        RAM[323] = 23'h672bc2;
        RAM[324] = 23'h674f2f;
        RAM[325] = 23'h677297;
        RAM[326] = 23'h6795fa;
        RAM[327] = 23'h67b957;
        RAM[328] = 23'h67dcae;
        RAM[329] = 23'h680000;
        RAM[330] = 23'h68234d;
        RAM[331] = 23'h684694;
        RAM[332] = 23'h6869d6;
        RAM[333] = 23'h688d13;
        RAM[334] = 23'h68b04a;
        RAM[335] = 23'h68d37c;
        RAM[336] = 23'h68f6a9;
        RAM[337] = 23'h6919d1;
        RAM[338] = 23'h693cf2;
        RAM[339] = 23'h69600f;
        RAM[340] = 23'h698327;
        RAM[341] = 23'h69a639;
        RAM[342] = 23'h69c946;
        RAM[343] = 23'h69ec4e;
        RAM[344] = 23'h6a0f50;
        RAM[345] = 23'h6a324e;
        RAM[346] = 23'h6a5546;
        RAM[347] = 23'h6a7839;
        RAM[348] = 23'h6a9b26;
        RAM[349] = 23'h6abe0f;
        RAM[350] = 23'h6ae0f2;
        RAM[351] = 23'h6b03d0;
        RAM[352] = 23'h6b26a9;
        RAM[353] = 23'h6b497d;
        RAM[354] = 23'h6b6c4b;
        RAM[355] = 23'h6b8f14;
        RAM[356] = 23'h6bb1d9;
        RAM[357] = 23'h6bd498;
        RAM[358] = 23'h6bf752;
        RAM[359] = 23'h6c1a07;
        RAM[360] = 23'h6c3cb7;
        RAM[361] = 23'h6c5f62;
        RAM[362] = 23'h6c8208;
        RAM[363] = 23'h6ca4a8;
        RAM[364] = 23'h6cc743;
        RAM[365] = 23'h6ce9da;
        RAM[366] = 23'h6d0c6c;
        RAM[367] = 23'h6d2ef8;
        RAM[368] = 23'h6d5180;
        RAM[369] = 23'h6d7402;
        RAM[370] = 23'h6d967f;
        RAM[371] = 23'h6db8f8;
        RAM[372] = 23'h6ddb6b;
        RAM[373] = 23'h6dfdd9;
        RAM[374] = 23'h6e2042;
        RAM[375] = 23'h6e42a7;
        RAM[376] = 23'h6e6507;
        RAM[377] = 23'h6e8761;
        RAM[378] = 23'h6ea9b6;
        RAM[379] = 23'h6ecc07;
        RAM[380] = 23'h6eee53;
        RAM[381] = 23'h6f1099;
        RAM[382] = 23'h6f32dc;
        RAM[383] = 23'h6f5519;
        RAM[384] = 23'h6f7751;
        RAM[385] = 23'h6f9983;
        RAM[386] = 23'h6fbbb2;
        RAM[387] = 23'h6fdddc;
        RAM[388] = 23'h700000;
        RAM[389] = 23'h702220;
        RAM[390] = 23'h70443b;
        RAM[391] = 23'h706651;
        RAM[392] = 23'h708862;
        RAM[393] = 23'h70aa6e;
        RAM[394] = 23'h70cc75;
        RAM[395] = 23'h70ee78;
        RAM[396] = 23'h711076;
        RAM[397] = 23'h713270;
        RAM[398] = 23'h715464;
        RAM[399] = 23'h717653;
        RAM[400] = 23'h71983e;
        RAM[401] = 23'h71ba24;
        RAM[402] = 23'h71dc06;
        RAM[403] = 23'h71fde2;
        RAM[404] = 23'h721fba;
        RAM[405] = 23'h72418d;
        RAM[406] = 23'h72635c;
        RAM[407] = 23'h728526;
        RAM[408] = 23'h72a6ea;
        RAM[409] = 23'h72c8ab;
        RAM[410] = 23'h72ea66;
        RAM[411] = 23'h730c1d;
        RAM[412] = 23'h732dd0;
        RAM[413] = 23'h734f7d;
        RAM[414] = 23'h737126;
        RAM[415] = 23'h7392ca;
        RAM[416] = 23'h73b46a;
        RAM[417] = 23'h73d605;
        RAM[418] = 23'h73f79b;
        RAM[419] = 23'h74192d;
        RAM[420] = 23'h743aba;
        RAM[421] = 23'h745c43;
        RAM[422] = 23'h747dc6;
        RAM[423] = 23'h749f45;
        RAM[424] = 23'h74c0c1;
        RAM[425] = 23'h74e237;
        RAM[426] = 23'h7503a8;
        RAM[427] = 23'h752515;
        RAM[428] = 23'h75467e;
        RAM[429] = 23'h7567e2;
        RAM[430] = 23'h758941;
        RAM[431] = 23'h75aa9b;
        RAM[432] = 23'h75cbf2;
        RAM[433] = 23'h75ed44;
        RAM[434] = 23'h760e91;
        RAM[435] = 23'h762fda;
        RAM[436] = 23'h76511e;
        RAM[437] = 23'h76725e;
        RAM[438] = 23'h76939a;
        RAM[439] = 23'h76b4d0;
        RAM[440] = 23'h76d603;
        RAM[441] = 23'h76f731;
        RAM[442] = 23'h77185a;
        RAM[443] = 23'h77397f;
        RAM[444] = 23'h775aa0;
        RAM[445] = 23'h777bbc;
        RAM[446] = 23'h779cd3;
        RAM[447] = 23'h77bde7;
        RAM[448] = 23'h77def5;
        RAM[449] = 23'h780000;
        RAM[450] = 23'h782106;
        RAM[451] = 23'h784208;
        RAM[452] = 23'h786305;
        RAM[453] = 23'h7883fe;
        RAM[454] = 23'h78a4f2;
        RAM[455] = 23'h78c5e3;
        RAM[456] = 23'h78e6ce;
        RAM[457] = 23'h7907b6;
        RAM[458] = 23'h792899;
        RAM[459] = 23'h794977;
        RAM[460] = 23'h796a52;
        RAM[461] = 23'h798b28;
        RAM[462] = 23'h79abfa;
        RAM[463] = 23'h79ccc8;
        RAM[464] = 23'h79ed91;
        RAM[465] = 23'h7a0e56;
        RAM[466] = 23'h7a2f16;
        RAM[467] = 23'h7a4fd3;
        RAM[468] = 23'h7a708b;
        RAM[469] = 23'h7a913e;
        RAM[470] = 23'h7ab1ee;
        RAM[471] = 23'h7ad299;
        RAM[472] = 23'h7af340;
        RAM[473] = 23'h7b13e3;
        RAM[474] = 23'h7b3481;
        RAM[475] = 23'h7b551b;
        RAM[476] = 23'h7b75b1;
        RAM[477] = 23'h7b9643;
        RAM[478] = 23'h7bb6d1;
        RAM[479] = 23'h7bd75a;
        RAM[480] = 23'h7bf7df;
        RAM[481] = 23'h7c1860;
        RAM[482] = 23'h7c38dd;
        RAM[483] = 23'h7c5956;
        RAM[484] = 23'h7c79ca;
        RAM[485] = 23'h7c9a3a;
        RAM[486] = 23'h7cbaa6;
        RAM[487] = 23'h7cdb0f;
        RAM[488] = 23'h7cfb72;
        RAM[489] = 23'h7d1bd2;
        RAM[490] = 23'h7d3c2d;
        RAM[491] = 23'h7d5c85;
        RAM[492] = 23'h7d7cd8;
        RAM[493] = 23'h7d9d27;
        RAM[494] = 23'h7dbd72;
        RAM[495] = 23'h7dddb9;
        RAM[496] = 23'h7dfdfc;
        RAM[497] = 23'h7e1e3b;
        RAM[498] = 23'h7e3e75;
        RAM[499] = 23'h7e5eab;
        RAM[500] = 23'h7e7ede;
        RAM[501] = 23'h7e9f0d;
        RAM[502] = 23'h7ebf37;
        RAM[503] = 23'h7edf5d;
        RAM[504] = 23'h7eff80;
        RAM[505] = 23'h7f1f9d;
        RAM[506] = 23'h7f3fb7;
        RAM[507] = 23'h7f5fcd;
        RAM[508] = 23'h7f7fdf;
        RAM[509] = 23'h7f9fed;
        RAM[510] = 23'h7fbff7;
        RAM[511] = 23'h7fdffd;
        RAM[512] = 23'h0;
        RAM[513] = 23'h1ffc;
        RAM[514] = 23'h3ff1;
        RAM[515] = 23'h5fdd;
        RAM[516] = 23'h7fc1;
        RAM[517] = 23'h9f9d;
        RAM[518] = 23'hbf71;
        RAM[519] = 23'hdf3e;
        RAM[520] = 23'hff02;
        RAM[521] = 23'h11ebf;
        RAM[522] = 23'h13e74;
        RAM[523] = 23'h15e22;
        RAM[524] = 23'h17dc7;
        RAM[525] = 23'h19d65;
        RAM[526] = 23'h1bcfb;
        RAM[527] = 23'h1dc89;
        RAM[528] = 23'h1fc10;
        RAM[529] = 23'h21b8f;
        RAM[530] = 23'h23b07;
        RAM[531] = 23'h25a77;
        RAM[532] = 23'h279de;
        RAM[533] = 23'h29940;
        RAM[534] = 23'h2b899;
        RAM[535] = 23'h2d7ea;
        RAM[536] = 23'h2f735;
        RAM[537] = 23'h31677;
        RAM[538] = 23'h335b3;
        RAM[539] = 23'h354e7;
        RAM[540] = 23'h37413;
        RAM[541] = 23'h39338;
        RAM[542] = 23'h3b256;
        RAM[543] = 23'h3d16d;
        RAM[544] = 23'h3f07b;
        RAM[545] = 23'h40f83;
        RAM[546] = 23'h42e84;
        RAM[547] = 23'h44d7d;
        RAM[548] = 23'h46c6f;
        RAM[549] = 23'h48b59;
        RAM[550] = 23'h4aa3d;
        RAM[551] = 23'h4c91a;
        RAM[552] = 23'h4e7ee;
        RAM[553] = 23'h506bd;
        RAM[554] = 23'h52583;
        RAM[555] = 23'h54444;
        RAM[556] = 23'h562fc;
        RAM[557] = 23'h581ad;
        RAM[558] = 23'h5a059;
        RAM[559] = 23'h5befc;
        RAM[560] = 23'h5dd98;
        RAM[561] = 23'h5fc2e;
        RAM[562] = 23'h61abd;
        RAM[563] = 23'h63944;
        RAM[564] = 23'h657c5;
        RAM[565] = 23'h6763f;
        RAM[566] = 23'h694b1;
        RAM[567] = 23'h6b31e;
        RAM[568] = 23'h6d183;
        RAM[569] = 23'h6efe1;
        RAM[570] = 23'h70e38;
        RAM[571] = 23'h72c89;
        RAM[572] = 23'h74ad3;
        RAM[573] = 23'h76916;
        RAM[574] = 23'h78752;
        RAM[575] = 23'h7a587;
        RAM[576] = 23'h7c3b7;
        RAM[577] = 23'h7e1df;
        RAM[578] = 23'h80000;
        RAM[579] = 23'h81e1b;
        RAM[580] = 23'h83c2f;
        RAM[581] = 23'h85a3d;
        RAM[582] = 23'h87844;
        RAM[583] = 23'h89644;
        RAM[584] = 23'h8b43e;
        RAM[585] = 23'h8d231;
        RAM[586] = 23'h8f01d;
        RAM[587] = 23'h90e03;
        RAM[588] = 23'h92be3;
        RAM[589] = 23'h949bb;
        RAM[590] = 23'h9678e;
        RAM[591] = 23'h9855a;
        RAM[592] = 23'h9a320;
        RAM[593] = 23'h9c0df;
        RAM[594] = 23'h9de98;
        RAM[595] = 23'h9fc4a;
        RAM[596] = 23'ha19f6;
        RAM[597] = 23'ha379c;
        RAM[598] = 23'ha553b;
        RAM[599] = 23'ha72d4;
        RAM[600] = 23'ha9066;
        RAM[601] = 23'haadf3;
        RAM[602] = 23'hacb79;
        RAM[603] = 23'hae8f9;
        RAM[604] = 23'hb0672;
        RAM[605] = 23'hb23e6;
        RAM[606] = 23'hb4153;
        RAM[607] = 23'hb5eb9;
        RAM[608] = 23'hb7c19;
        RAM[609] = 23'hb9974;
        RAM[610] = 23'hbb6c8;
        RAM[611] = 23'hbd417;
        RAM[612] = 23'hbf15e;
        RAM[613] = 23'hc0ea0;
        RAM[614] = 23'hc2bdc;
        RAM[615] = 23'hc4912;
        RAM[616] = 23'hc6641;
        RAM[617] = 23'hc836b;
        RAM[618] = 23'hca08e;
        RAM[619] = 23'hcbdab;
        RAM[620] = 23'hcdac3;
        RAM[621] = 23'hcf7d4;
        RAM[622] = 23'hd14e0;
        RAM[623] = 23'hd31e5;
        RAM[624] = 23'hd4ee4;
        RAM[625] = 23'hd6bde;
        RAM[626] = 23'hd88d2;
        RAM[627] = 23'hda5bf;
        RAM[628] = 23'hdc2a7;
        RAM[629] = 23'hddf89;
        RAM[630] = 23'hdfc65;
        RAM[631] = 23'he193b;
        RAM[632] = 23'he360c;
        RAM[633] = 23'he52d6;
        RAM[634] = 23'he6f9b;
        RAM[635] = 23'he8c5a;
        RAM[636] = 23'hea913;
        RAM[637] = 23'hec5c6;
        RAM[638] = 23'hee273;
        RAM[639] = 23'heff1b;
        RAM[640] = 23'hf1bbd;
        RAM[641] = 23'hf3859;
        RAM[642] = 23'hf54f0;
        RAM[643] = 23'hf7181;
        RAM[644] = 23'hf8e0c;
        RAM[645] = 23'hfaa91;
        RAM[646] = 23'hfc711;
        RAM[647] = 23'hfe38c;
        RAM[648] = 23'h100000;
        RAM[649] = 23'h101c6f;
        RAM[650] = 23'h1038d9;
        RAM[651] = 23'h10553c;
        RAM[652] = 23'h10719a;
        RAM[653] = 23'h108df3;
        RAM[654] = 23'h10aa46;
        RAM[655] = 23'h10c694;
        RAM[656] = 23'h10e2db;
        RAM[657] = 23'h10ff1e;
        RAM[658] = 23'h111b5b;
        RAM[659] = 23'h113792;
        RAM[660] = 23'h1153c5;
        RAM[661] = 23'h116ff1;
        RAM[662] = 23'h118c18;
        RAM[663] = 23'h11a83a;
        RAM[664] = 23'h11c456;
        RAM[665] = 23'h11e06d;
        RAM[666] = 23'h11fc7e;
        RAM[667] = 23'h12188a;
        RAM[668] = 23'h123491;
        RAM[669] = 23'h125092;
        RAM[670] = 23'h126c8e;
        RAM[671] = 23'h128885;
        RAM[672] = 23'h12a476;
        RAM[673] = 23'h12c061;
        RAM[674] = 23'h12dc48;
        RAM[675] = 23'h12f82a;
        RAM[676] = 23'h131405;
        RAM[677] = 23'h132fdc;
        RAM[678] = 23'h134bae;
        RAM[679] = 23'h13677a;
        RAM[680] = 23'h138341;
        RAM[681] = 23'h139f02;
        RAM[682] = 23'h13babf;
        RAM[683] = 23'h13d677;
        RAM[684] = 23'h13f229;
        RAM[685] = 23'h140dd6;
        RAM[686] = 23'h14297d;
        RAM[687] = 23'h144520;
        RAM[688] = 23'h1460be;
        RAM[689] = 23'h147c56;
        RAM[690] = 23'h1497ea;
        RAM[691] = 23'h14b378;
        RAM[692] = 23'h14cf01;
        RAM[693] = 23'h14ea85;
        RAM[694] = 23'h150603;
        RAM[695] = 23'h15217d;
        RAM[696] = 23'h153cf2;
        RAM[697] = 23'h155862;
        RAM[698] = 23'h1573cc;
        RAM[699] = 23'h158f32;
        RAM[700] = 23'h15aa92;
        RAM[701] = 23'h15c5ee;
        RAM[702] = 23'h15e145;
        RAM[703] = 23'h15fc96;
        RAM[704] = 23'h1617e3;
        RAM[705] = 23'h16332b;
        RAM[706] = 23'h164e6d;
        RAM[707] = 23'h1669ab;
        RAM[708] = 23'h1684e4;
        RAM[709] = 23'h16a018;
        RAM[710] = 23'h16bb47;
        RAM[711] = 23'h16d671;
        RAM[712] = 23'h16f196;
        RAM[713] = 23'h170cb7;
        RAM[714] = 23'h1727d2;
        RAM[715] = 23'h1742e9;
        RAM[716] = 23'h175dfb;
        RAM[717] = 23'h177908;
        RAM[718] = 23'h179410;
        RAM[719] = 23'h17af13;
        RAM[720] = 23'h17ca11;
        RAM[721] = 23'h17e50b;
        RAM[722] = 23'h180000;
        RAM[723] = 23'h181af0;
        RAM[724] = 23'h1835db;
        RAM[725] = 23'h1850c2;
        RAM[726] = 23'h186ba4;
        RAM[727] = 23'h188681;
        RAM[728] = 23'h18a15a;
        RAM[729] = 23'h18bc2d;
        RAM[730] = 23'h18d6fc;
        RAM[731] = 23'h18f1c6;
        RAM[732] = 23'h190c8c;
        RAM[733] = 23'h19274d;
        RAM[734] = 23'h194209;
        RAM[735] = 23'h195cc1;
        RAM[736] = 23'h197773;
        RAM[737] = 23'h199222;
        RAM[738] = 23'h19accc;
        RAM[739] = 23'h19c770;
        RAM[740] = 23'h19e211;
        RAM[741] = 23'h19fcad;
        RAM[742] = 23'h1a1744;
        RAM[743] = 23'h1a31d7;
        RAM[744] = 23'h1a4c65;
        RAM[745] = 23'h1a66ee;
        RAM[746] = 23'h1a8173;
        RAM[747] = 23'h1a9bf4;
        RAM[748] = 23'h1ab66f;
        RAM[749] = 23'h1ad0e7;
        RAM[750] = 23'h1aeb5a;
        RAM[751] = 23'h1b05c7;
        RAM[752] = 23'h1b2032;
        RAM[753] = 23'h1b3a97;
        RAM[754] = 23'h1b54f8;
        RAM[755] = 23'h1b6f54;
        RAM[756] = 23'h1b89ac;
        RAM[757] = 23'h1ba3ff;
        RAM[758] = 23'h1bbe4e;
        RAM[759] = 23'h1bd899;
        RAM[760] = 23'h1bf2df;
        RAM[761] = 23'h1c0d20;
        RAM[762] = 23'h1c275e;
        RAM[763] = 23'h1c4196;
        RAM[764] = 23'h1c5bca;
        RAM[765] = 23'h1c75fb;
        RAM[766] = 23'h1c9026;
        RAM[767] = 23'h1caa4e;
        RAM[768] = 23'h1cc471;
        RAM[769] = 23'h1cde8f;
        RAM[770] = 23'h1cf8a9;
        RAM[771] = 23'h1d12bf;
        RAM[772] = 23'h1d2cd1;
        RAM[773] = 23'h1d46de;
        RAM[774] = 23'h1d60e7;
        RAM[775] = 23'h1d7aec;
        RAM[776] = 23'h1d94ec;
        RAM[777] = 23'h1daee8;
        RAM[778] = 23'h1dc8e0;
        RAM[779] = 23'h1de2d3;
        RAM[780] = 23'h1dfcc2;
        RAM[781] = 23'h1e16ad;
        RAM[782] = 23'h1e3094;
        RAM[783] = 23'h1e4a77;
        RAM[784] = 23'h1e6455;
        RAM[785] = 23'h1e7e2f;
        RAM[786] = 23'h1e9805;
        RAM[787] = 23'h1eb1d6;
        RAM[788] = 23'h1ecba4;
        RAM[789] = 23'h1ee56d;
        RAM[790] = 23'h1eff32;
        RAM[791] = 23'h1f18f2;
        RAM[792] = 23'h1f32af;
        RAM[793] = 23'h1f4c68;
        RAM[794] = 23'h1f661c;
        RAM[795] = 23'h1f7fcc;
        RAM[796] = 23'h1f9978;
        RAM[797] = 23'h1fb320;
        RAM[798] = 23'h1fccc5;
        RAM[799] = 23'h1fe664;
        RAM[800] = 23'h200000;
        RAM[801] = 23'h201998;
        RAM[802] = 23'h20332b;
        RAM[803] = 23'h204cba;
        RAM[804] = 23'h206646;
        RAM[805] = 23'h207fcd;
        RAM[806] = 23'h209950;
        RAM[807] = 23'h20b2cf;
        RAM[808] = 23'h20cc4a;
        RAM[809] = 23'h20e5c1;
        RAM[810] = 23'h20ff34;
        RAM[811] = 23'h2118a3;
        RAM[812] = 23'h21320e;
        RAM[813] = 23'h214b75;
        RAM[814] = 23'h2164d8;
        RAM[815] = 23'h217e37;
        RAM[816] = 23'h219792;
        RAM[817] = 23'h21b0ea;
        RAM[818] = 23'h21ca3d;
        RAM[819] = 23'h21e38c;
        RAM[820] = 23'h21fcd7;
        RAM[821] = 23'h22161e;
        RAM[822] = 23'h222f61;
        RAM[823] = 23'h2248a1;
        RAM[824] = 23'h2261dc;
        RAM[825] = 23'h227b14;
        RAM[826] = 23'h229447;
        RAM[827] = 23'h22ad76;
        RAM[828] = 23'h22c6a2;
        RAM[829] = 23'h22dfca;
        RAM[830] = 23'h22f8ee;
        RAM[831] = 23'h23120e;
        RAM[832] = 23'h232b2a;
        RAM[833] = 23'h234443;
        RAM[834] = 23'h235d58;
        RAM[835] = 23'h237668;
        RAM[836] = 23'h238f75;
        RAM[837] = 23'h23a87e;
        RAM[838] = 23'h23c184;
        RAM[839] = 23'h23da85;
        RAM[840] = 23'h23f383;
        RAM[841] = 23'h240c7c;
        RAM[842] = 23'h242572;
        RAM[843] = 23'h243e64;
        RAM[844] = 23'h245753;
        RAM[845] = 23'h24703d;
        RAM[846] = 23'h248924;
        RAM[847] = 23'h24a207;
        RAM[848] = 23'h24bae7;
        RAM[849] = 23'h24d3c2;
        RAM[850] = 23'h24ec9a;
        RAM[851] = 23'h25056e;
        RAM[852] = 23'h251e3e;
        RAM[853] = 23'h25370b;
        RAM[854] = 23'h254fd4;
        RAM[855] = 23'h256899;
        RAM[856] = 23'h25815a;
        RAM[857] = 23'h259a18;
        RAM[858] = 23'h25b2d2;
        RAM[859] = 23'h25cb89;
        RAM[860] = 23'h25e43b;
        RAM[861] = 23'h25fcea;
        RAM[862] = 23'h261596;
        RAM[863] = 23'h262e3d;
        RAM[864] = 23'h2646e1;
        RAM[865] = 23'h265f82;
        RAM[866] = 23'h26781f;
        RAM[867] = 23'h2690b8;
        RAM[868] = 23'h26a94d;
        RAM[869] = 23'h26c1df;
        RAM[870] = 23'h26da6d;
        RAM[871] = 23'h26f2f8;
        RAM[872] = 23'h270b7f;
        RAM[873] = 23'h272402;
        RAM[874] = 23'h273c82;
        RAM[875] = 23'h2754fe;
        RAM[876] = 23'h276d77;
        RAM[877] = 23'h2785eb;
        RAM[878] = 23'h279e5d;
        RAM[879] = 23'h27b6cb;
        RAM[880] = 23'h27cf36;
        RAM[881] = 23'h27e79d;
        RAM[882] = 23'h280000;
        RAM[883] = 23'h281860;
        RAM[884] = 23'h2830bc;
        RAM[885] = 23'h284915;
        RAM[886] = 23'h286169;
        RAM[887] = 23'h2879bb;
        RAM[888] = 23'h289209;
        RAM[889] = 23'h28aa54;
        RAM[890] = 23'h28c29b;
        RAM[891] = 23'h28dadf;
        RAM[892] = 23'h28f31f;
        RAM[893] = 23'h290b5c;
        RAM[894] = 23'h292395;
        RAM[895] = 23'h293bcb;
        RAM[896] = 23'h2953fd;
        RAM[897] = 23'h296c2c;
        RAM[898] = 23'h298457;
        RAM[899] = 23'h299c7f;
        RAM[900] = 23'h29b4a4;
        RAM[901] = 23'h29ccc5;
        RAM[902] = 23'h29e4e3;
        RAM[903] = 23'h29fcfd;
        RAM[904] = 23'h2a1514;
        RAM[905] = 23'h2a2d27;
        RAM[906] = 23'h2a4537;
        RAM[907] = 23'h2a5d44;
        RAM[908] = 23'h2a754d;
        RAM[909] = 23'h2a8d53;
        RAM[910] = 23'h2aa555;
        RAM[911] = 23'h2abd54;
        RAM[912] = 23'h2ad550;
        RAM[913] = 23'h2aed48;
        RAM[914] = 23'h2b053d;
        RAM[915] = 23'h2b1d2f;
        RAM[916] = 23'h2b351d;
        RAM[917] = 23'h2b4d08;
        RAM[918] = 23'h2b64f0;
        RAM[919] = 23'h2b7cd4;
        RAM[920] = 23'h2b94b5;
        RAM[921] = 23'h2bac92;
        RAM[922] = 23'h2bc46d;
        RAM[923] = 23'h2bdc44;
        RAM[924] = 23'h2bf417;
        RAM[925] = 23'h2c0be8;
        RAM[926] = 23'h2c23b5;
        RAM[927] = 23'h2c3b7f;
        RAM[928] = 23'h2c5345;
        RAM[929] = 23'h2c6b08;
        RAM[930] = 23'h2c82c8;
        RAM[931] = 23'h2c9a85;
        RAM[932] = 23'h2cb23e;
        RAM[933] = 23'h2cc9f5;
        RAM[934] = 23'h2ce1a7;
        RAM[935] = 23'h2cf957;
        RAM[936] = 23'h2d1104;
        RAM[937] = 23'h2d28ad;
        RAM[938] = 23'h2d4053;
        RAM[939] = 23'h2d57f5;
        RAM[940] = 23'h2d6f94;
        RAM[941] = 23'h2d8731;
        RAM[942] = 23'h2d9eca;
        RAM[943] = 23'h2db660;
        RAM[944] = 23'h2dcdf3;
        RAM[945] = 23'h2de582;
        RAM[946] = 23'h2dfd0f;
        RAM[947] = 23'h2e1497;
        RAM[948] = 23'h2e2c1d;
        RAM[949] = 23'h2e43a0;
        RAM[950] = 23'h2e5b20;
        RAM[951] = 23'h2e729c;
        RAM[952] = 23'h2e8a15;
        RAM[953] = 23'h2ea18c;
        RAM[954] = 23'h2eb8fe;
        RAM[955] = 23'h2ed06e;
        RAM[956] = 23'h2ee7db;
        RAM[957] = 23'h2eff45;
        RAM[958] = 23'h2f16ab;
        RAM[959] = 23'h2f2e0e;
        RAM[960] = 23'h2f456e;
        RAM[961] = 23'h2f5ccb;
        RAM[962] = 23'h2f7425;
        RAM[963] = 23'h2f8b7c;
        RAM[964] = 23'h2fa2d0;
        RAM[965] = 23'h2fba21;
        RAM[966] = 23'h2fd16e;
        RAM[967] = 23'h2fe8b9;
        RAM[968] = 23'h300000;
        RAM[969] = 23'h301744;
        RAM[970] = 23'h302e85;
        RAM[971] = 23'h3045c4;
        RAM[972] = 23'h305cfe;
        RAM[973] = 23'h307437;
        RAM[974] = 23'h308b6b;
        RAM[975] = 23'h30a29d;
        RAM[976] = 23'h30b9cc;
        RAM[977] = 23'h30d0f8;
        RAM[978] = 23'h30e821;
        RAM[979] = 23'h30ff47;
        RAM[980] = 23'h311669;
        RAM[981] = 23'h312d89;
        RAM[982] = 23'h3144a5;
        RAM[983] = 23'h315bbf;
        RAM[984] = 23'h3172d6;
        RAM[985] = 23'h3189ea;
        RAM[986] = 23'h31a0fb;
        RAM[987] = 23'h31b808;
        RAM[988] = 23'h31cf13;
        RAM[989] = 23'h31e61b;
        RAM[990] = 23'h31fd1f;
        RAM[991] = 23'h321421;
        RAM[992] = 23'h322b20;
        RAM[993] = 23'h32421c;
        RAM[994] = 23'h325915;
        RAM[995] = 23'h32700b;
        RAM[996] = 23'h3286fe;
        RAM[997] = 23'h329dee;
        RAM[998] = 23'h32b4db;
        RAM[999] = 23'h32cbc5;
        RAM[1000] = 23'h32e2ac;
        RAM[1001] = 23'h32f990;
        RAM[1002] = 23'h331071;
        RAM[1003] = 23'h332750;
        RAM[1004] = 23'h333e2b;
        RAM[1005] = 23'h335503;
        RAM[1006] = 23'h336bda;
        RAM[1007] = 23'h3382ac;
        RAM[1008] = 23'h33997c;
        RAM[1009] = 23'h33b049;
        RAM[1010] = 23'h33c713;
        RAM[1011] = 23'h33ddda;
        RAM[1012] = 23'h33f49f;
        RAM[1013] = 23'h340b60;
        RAM[1014] = 23'h34221e;
        RAM[1015] = 23'h3438da;
        RAM[1016] = 23'h344f93;
        RAM[1017] = 23'h346649;
        RAM[1018] = 23'h347cfc;
        RAM[1019] = 23'h3493ad;
        RAM[1020] = 23'h34aa5a;
        RAM[1021] = 23'h34c104;
        RAM[1022] = 23'h34d7ac;
        RAM[1023] = 23'h34ee51;
    end
endmodule

module fsqrt_grad_table (
    input wire clk, 
    input wire [9:0] addr,
    output reg [12:0] grd);

    reg [12:0] RAM [1023:0];
    always @(posedge clk)
        grd <= RAM[addr];
    initial begin
        RAM[0] = 13'h169d;
        RAM[1] = 13'h1698;
        RAM[2] = 13'h1692;
        RAM[3] = 13'h168c;
        RAM[4] = 13'h1687;
        RAM[5] = 13'h1681;
        RAM[6] = 13'h167c;
        RAM[7] = 13'h1676;
        RAM[8] = 13'h1671;
        RAM[9] = 13'h166b;
        RAM[10] = 13'h1666;
        RAM[11] = 13'h1660;
        RAM[12] = 13'h165b;
        RAM[13] = 13'h1655;
        RAM[14] = 13'h1650;
        RAM[15] = 13'h164a;
        RAM[16] = 13'h1645;
        RAM[17] = 13'h1640;
        RAM[18] = 13'h163a;
        RAM[19] = 13'h1635;
        RAM[20] = 13'h1630;
        RAM[21] = 13'h162a;
        RAM[22] = 13'h1625;
        RAM[23] = 13'h1620;
        RAM[24] = 13'h161a;
        RAM[25] = 13'h1615;
        RAM[26] = 13'h1610;
        RAM[27] = 13'h160b;
        RAM[28] = 13'h1605;
        RAM[29] = 13'h1600;
        RAM[30] = 13'h15fb;
        RAM[31] = 13'h15f6;
        RAM[32] = 13'h15f1;
        RAM[33] = 13'h15eb;
        RAM[34] = 13'h15e6;
        RAM[35] = 13'h15e1;
        RAM[36] = 13'h15dc;
        RAM[37] = 13'h15d7;
        RAM[38] = 13'h15d2;
        RAM[39] = 13'h15cd;
        RAM[40] = 13'h15c8;
        RAM[41] = 13'h15c3;
        RAM[42] = 13'h15be;
        RAM[43] = 13'h15b9;
        RAM[44] = 13'h15b4;
        RAM[45] = 13'h15af;
        RAM[46] = 13'h15aa;
        RAM[47] = 13'h15a5;
        RAM[48] = 13'h15a0;
        RAM[49] = 13'h159b;
        RAM[50] = 13'h1596;
        RAM[51] = 13'h1591;
        RAM[52] = 13'h158c;
        RAM[53] = 13'h1587;
        RAM[54] = 13'h1582;
        RAM[55] = 13'h157e;
        RAM[56] = 13'h1579;
        RAM[57] = 13'h1574;
        RAM[58] = 13'h156f;
        RAM[59] = 13'h156a;
        RAM[60] = 13'h1566;
        RAM[61] = 13'h1561;
        RAM[62] = 13'h155c;
        RAM[63] = 13'h1557;
        RAM[64] = 13'h1552;
        RAM[65] = 13'h154e;
        RAM[66] = 13'h1549;
        RAM[67] = 13'h1544;
        RAM[68] = 13'h1540;
        RAM[69] = 13'h153b;
        RAM[70] = 13'h1536;
        RAM[71] = 13'h1532;
        RAM[72] = 13'h152d;
        RAM[73] = 13'h1528;
        RAM[74] = 13'h1524;
        RAM[75] = 13'h151f;
        RAM[76] = 13'h151b;
        RAM[77] = 13'h1516;
        RAM[78] = 13'h1511;
        RAM[79] = 13'h150d;
        RAM[80] = 13'h1508;
        RAM[81] = 13'h1504;
        RAM[82] = 13'h14ff;
        RAM[83] = 13'h14fb;
        RAM[84] = 13'h14f6;
        RAM[85] = 13'h14f2;
        RAM[86] = 13'h14ed;
        RAM[87] = 13'h14e9;
        RAM[88] = 13'h14e4;
        RAM[89] = 13'h14e0;
        RAM[90] = 13'h14db;
        RAM[91] = 13'h14d7;
        RAM[92] = 13'h14d3;
        RAM[93] = 13'h14ce;
        RAM[94] = 13'h14ca;
        RAM[95] = 13'h14c5;
        RAM[96] = 13'h14c1;
        RAM[97] = 13'h14bd;
        RAM[98] = 13'h14b8;
        RAM[99] = 13'h14b4;
        RAM[100] = 13'h14b0;
        RAM[101] = 13'h14ab;
        RAM[102] = 13'h14a7;
        RAM[103] = 13'h14a3;
        RAM[104] = 13'h149e;
        RAM[105] = 13'h149a;
        RAM[106] = 13'h1496;
        RAM[107] = 13'h1492;
        RAM[108] = 13'h148d;
        RAM[109] = 13'h1489;
        RAM[110] = 13'h1485;
        RAM[111] = 13'h1481;
        RAM[112] = 13'h147c;
        RAM[113] = 13'h1478;
        RAM[114] = 13'h1474;
        RAM[115] = 13'h1470;
        RAM[116] = 13'h146c;
        RAM[117] = 13'h1468;
        RAM[118] = 13'h1463;
        RAM[119] = 13'h145f;
        RAM[120] = 13'h145b;
        RAM[121] = 13'h1457;
        RAM[122] = 13'h1453;
        RAM[123] = 13'h144f;
        RAM[124] = 13'h144b;
        RAM[125] = 13'h1447;
        RAM[126] = 13'h1443;
        RAM[127] = 13'h143f;
        RAM[128] = 13'h143b;
        RAM[129] = 13'h1437;
        RAM[130] = 13'h1432;
        RAM[131] = 13'h142e;
        RAM[132] = 13'h142a;
        RAM[133] = 13'h1426;
        RAM[134] = 13'h1422;
        RAM[135] = 13'h141e;
        RAM[136] = 13'h141b;
        RAM[137] = 13'h1417;
        RAM[138] = 13'h1413;
        RAM[139] = 13'h140f;
        RAM[140] = 13'h140b;
        RAM[141] = 13'h1407;
        RAM[142] = 13'h1403;
        RAM[143] = 13'h13ff;
        RAM[144] = 13'h13fb;
        RAM[145] = 13'h13f7;
        RAM[146] = 13'h13f3;
        RAM[147] = 13'h13ef;
        RAM[148] = 13'h13ec;
        RAM[149] = 13'h13e8;
        RAM[150] = 13'h13e4;
        RAM[151] = 13'h13e0;
        RAM[152] = 13'h13dc;
        RAM[153] = 13'h13d8;
        RAM[154] = 13'h13d5;
        RAM[155] = 13'h13d1;
        RAM[156] = 13'h13cd;
        RAM[157] = 13'h13c9;
        RAM[158] = 13'h13c5;
        RAM[159] = 13'h13c2;
        RAM[160] = 13'h13be;
        RAM[161] = 13'h13ba;
        RAM[162] = 13'h13b6;
        RAM[163] = 13'h13b3;
        RAM[164] = 13'h13af;
        RAM[165] = 13'h13ab;
        RAM[166] = 13'h13a7;
        RAM[167] = 13'h13a4;
        RAM[168] = 13'h13a0;
        RAM[169] = 13'h139c;
        RAM[170] = 13'h1399;
        RAM[171] = 13'h1395;
        RAM[172] = 13'h1391;
        RAM[173] = 13'h138e;
        RAM[174] = 13'h138a;
        RAM[175] = 13'h1386;
        RAM[176] = 13'h1383;
        RAM[177] = 13'h137f;
        RAM[178] = 13'h137c;
        RAM[179] = 13'h1378;
        RAM[180] = 13'h1374;
        RAM[181] = 13'h1371;
        RAM[182] = 13'h136d;
        RAM[183] = 13'h136a;
        RAM[184] = 13'h1366;
        RAM[185] = 13'h1362;
        RAM[186] = 13'h135f;
        RAM[187] = 13'h135b;
        RAM[188] = 13'h1358;
        RAM[189] = 13'h1354;
        RAM[190] = 13'h1351;
        RAM[191] = 13'h134d;
        RAM[192] = 13'h134a;
        RAM[193] = 13'h1346;
        RAM[194] = 13'h1343;
        RAM[195] = 13'h133f;
        RAM[196] = 13'h133c;
        RAM[197] = 13'h1338;
        RAM[198] = 13'h1335;
        RAM[199] = 13'h1331;
        RAM[200] = 13'h132e;
        RAM[201] = 13'h132a;
        RAM[202] = 13'h1327;
        RAM[203] = 13'h1324;
        RAM[204] = 13'h1320;
        RAM[205] = 13'h131d;
        RAM[206] = 13'h1319;
        RAM[207] = 13'h1316;
        RAM[208] = 13'h1313;
        RAM[209] = 13'h130f;
        RAM[210] = 13'h130c;
        RAM[211] = 13'h1308;
        RAM[212] = 13'h1305;
        RAM[213] = 13'h1302;
        RAM[214] = 13'h12fe;
        RAM[215] = 13'h12fb;
        RAM[216] = 13'h12f8;
        RAM[217] = 13'h12f4;
        RAM[218] = 13'h12f1;
        RAM[219] = 13'h12ee;
        RAM[220] = 13'h12ea;
        RAM[221] = 13'h12e7;
        RAM[222] = 13'h12e4;
        RAM[223] = 13'h12e1;
        RAM[224] = 13'h12dd;
        RAM[225] = 13'h12da;
        RAM[226] = 13'h12d7;
        RAM[227] = 13'h12d3;
        RAM[228] = 13'h12d0;
        RAM[229] = 13'h12cd;
        RAM[230] = 13'h12ca;
        RAM[231] = 13'h12c6;
        RAM[232] = 13'h12c3;
        RAM[233] = 13'h12c0;
        RAM[234] = 13'h12bd;
        RAM[235] = 13'h12ba;
        RAM[236] = 13'h12b6;
        RAM[237] = 13'h12b3;
        RAM[238] = 13'h12b0;
        RAM[239] = 13'h12ad;
        RAM[240] = 13'h12aa;
        RAM[241] = 13'h12a6;
        RAM[242] = 13'h12a3;
        RAM[243] = 13'h12a0;
        RAM[244] = 13'h129d;
        RAM[245] = 13'h129a;
        RAM[246] = 13'h1297;
        RAM[247] = 13'h1294;
        RAM[248] = 13'h1290;
        RAM[249] = 13'h128d;
        RAM[250] = 13'h128a;
        RAM[251] = 13'h1287;
        RAM[252] = 13'h1284;
        RAM[253] = 13'h1281;
        RAM[254] = 13'h127e;
        RAM[255] = 13'h127b;
        RAM[256] = 13'h1278;
        RAM[257] = 13'h1275;
        RAM[258] = 13'h1271;
        RAM[259] = 13'h126e;
        RAM[260] = 13'h126b;
        RAM[261] = 13'h1268;
        RAM[262] = 13'h1265;
        RAM[263] = 13'h1262;
        RAM[264] = 13'h125f;
        RAM[265] = 13'h125c;
        RAM[266] = 13'h1259;
        RAM[267] = 13'h1256;
        RAM[268] = 13'h1253;
        RAM[269] = 13'h1250;
        RAM[270] = 13'h124d;
        RAM[271] = 13'h124a;
        RAM[272] = 13'h1247;
        RAM[273] = 13'h1244;
        RAM[274] = 13'h1241;
        RAM[275] = 13'h123e;
        RAM[276] = 13'h123b;
        RAM[277] = 13'h1238;
        RAM[278] = 13'h1235;
        RAM[279] = 13'h1232;
        RAM[280] = 13'h122f;
        RAM[281] = 13'h122d;
        RAM[282] = 13'h122a;
        RAM[283] = 13'h1227;
        RAM[284] = 13'h1224;
        RAM[285] = 13'h1221;
        RAM[286] = 13'h121e;
        RAM[287] = 13'h121b;
        RAM[288] = 13'h1218;
        RAM[289] = 13'h1215;
        RAM[290] = 13'h1212;
        RAM[291] = 13'h120f;
        RAM[292] = 13'h120d;
        RAM[293] = 13'h120a;
        RAM[294] = 13'h1207;
        RAM[295] = 13'h1204;
        RAM[296] = 13'h1201;
        RAM[297] = 13'h11fe;
        RAM[298] = 13'h11fb;
        RAM[299] = 13'h11f9;
        RAM[300] = 13'h11f6;
        RAM[301] = 13'h11f3;
        RAM[302] = 13'h11f0;
        RAM[303] = 13'h11ed;
        RAM[304] = 13'h11eb;
        RAM[305] = 13'h11e8;
        RAM[306] = 13'h11e5;
        RAM[307] = 13'h11e2;
        RAM[308] = 13'h11df;
        RAM[309] = 13'h11dd;
        RAM[310] = 13'h11da;
        RAM[311] = 13'h11d7;
        RAM[312] = 13'h11d4;
        RAM[313] = 13'h11d1;
        RAM[314] = 13'h11cf;
        RAM[315] = 13'h11cc;
        RAM[316] = 13'h11c9;
        RAM[317] = 13'h11c6;
        RAM[318] = 13'h11c4;
        RAM[319] = 13'h11c1;
        RAM[320] = 13'h11be;
        RAM[321] = 13'h11bc;
        RAM[322] = 13'h11b9;
        RAM[323] = 13'h11b6;
        RAM[324] = 13'h11b3;
        RAM[325] = 13'h11b1;
        RAM[326] = 13'h11ae;
        RAM[327] = 13'h11ab;
        RAM[328] = 13'h11a9;
        RAM[329] = 13'h11a6;
        RAM[330] = 13'h11a3;
        RAM[331] = 13'h11a1;
        RAM[332] = 13'h119e;
        RAM[333] = 13'h119b;
        RAM[334] = 13'h1199;
        RAM[335] = 13'h1196;
        RAM[336] = 13'h1193;
        RAM[337] = 13'h1191;
        RAM[338] = 13'h118e;
        RAM[339] = 13'h118b;
        RAM[340] = 13'h1189;
        RAM[341] = 13'h1186;
        RAM[342] = 13'h1183;
        RAM[343] = 13'h1181;
        RAM[344] = 13'h117e;
        RAM[345] = 13'h117c;
        RAM[346] = 13'h1179;
        RAM[347] = 13'h1176;
        RAM[348] = 13'h1174;
        RAM[349] = 13'h1171;
        RAM[350] = 13'h116f;
        RAM[351] = 13'h116c;
        RAM[352] = 13'h1169;
        RAM[353] = 13'h1167;
        RAM[354] = 13'h1164;
        RAM[355] = 13'h1162;
        RAM[356] = 13'h115f;
        RAM[357] = 13'h115d;
        RAM[358] = 13'h115a;
        RAM[359] = 13'h1157;
        RAM[360] = 13'h1155;
        RAM[361] = 13'h1152;
        RAM[362] = 13'h1150;
        RAM[363] = 13'h114d;
        RAM[364] = 13'h114b;
        RAM[365] = 13'h1148;
        RAM[366] = 13'h1146;
        RAM[367] = 13'h1143;
        RAM[368] = 13'h1141;
        RAM[369] = 13'h113e;
        RAM[370] = 13'h113c;
        RAM[371] = 13'h1139;
        RAM[372] = 13'h1137;
        RAM[373] = 13'h1134;
        RAM[374] = 13'h1132;
        RAM[375] = 13'h112f;
        RAM[376] = 13'h112d;
        RAM[377] = 13'h112a;
        RAM[378] = 13'h1128;
        RAM[379] = 13'h1125;
        RAM[380] = 13'h1123;
        RAM[381] = 13'h1120;
        RAM[382] = 13'h111e;
        RAM[383] = 13'h111c;
        RAM[384] = 13'h1119;
        RAM[385] = 13'h1117;
        RAM[386] = 13'h1114;
        RAM[387] = 13'h1112;
        RAM[388] = 13'h110f;
        RAM[389] = 13'h110d;
        RAM[390] = 13'h110b;
        RAM[391] = 13'h1108;
        RAM[392] = 13'h1106;
        RAM[393] = 13'h1103;
        RAM[394] = 13'h1101;
        RAM[395] = 13'h10fe;
        RAM[396] = 13'h10fc;
        RAM[397] = 13'h10fa;
        RAM[398] = 13'h10f7;
        RAM[399] = 13'h10f5;
        RAM[400] = 13'h10f3;
        RAM[401] = 13'h10f0;
        RAM[402] = 13'h10ee;
        RAM[403] = 13'h10eb;
        RAM[404] = 13'h10e9;
        RAM[405] = 13'h10e7;
        RAM[406] = 13'h10e4;
        RAM[407] = 13'h10e2;
        RAM[408] = 13'h10e0;
        RAM[409] = 13'h10dd;
        RAM[410] = 13'h10db;
        RAM[411] = 13'h10d9;
        RAM[412] = 13'h10d6;
        RAM[413] = 13'h10d4;
        RAM[414] = 13'h10d2;
        RAM[415] = 13'h10cf;
        RAM[416] = 13'h10cd;
        RAM[417] = 13'h10cb;
        RAM[418] = 13'h10c8;
        RAM[419] = 13'h10c6;
        RAM[420] = 13'h10c4;
        RAM[421] = 13'h10c1;
        RAM[422] = 13'h10bf;
        RAM[423] = 13'h10bd;
        RAM[424] = 13'h10bb;
        RAM[425] = 13'h10b8;
        RAM[426] = 13'h10b6;
        RAM[427] = 13'h10b4;
        RAM[428] = 13'h10b1;
        RAM[429] = 13'h10af;
        RAM[430] = 13'h10ad;
        RAM[431] = 13'h10ab;
        RAM[432] = 13'h10a8;
        RAM[433] = 13'h10a6;
        RAM[434] = 13'h10a4;
        RAM[435] = 13'h10a2;
        RAM[436] = 13'h109f;
        RAM[437] = 13'h109d;
        RAM[438] = 13'h109b;
        RAM[439] = 13'h1099;
        RAM[440] = 13'h1096;
        RAM[441] = 13'h1094;
        RAM[442] = 13'h1092;
        RAM[443] = 13'h1090;
        RAM[444] = 13'h108e;
        RAM[445] = 13'h108b;
        RAM[446] = 13'h1089;
        RAM[447] = 13'h1087;
        RAM[448] = 13'h1085;
        RAM[449] = 13'h1083;
        RAM[450] = 13'h1080;
        RAM[451] = 13'h107e;
        RAM[452] = 13'h107c;
        RAM[453] = 13'h107a;
        RAM[454] = 13'h1078;
        RAM[455] = 13'h1075;
        RAM[456] = 13'h1073;
        RAM[457] = 13'h1071;
        RAM[458] = 13'h106f;
        RAM[459] = 13'h106d;
        RAM[460] = 13'h106b;
        RAM[461] = 13'h1068;
        RAM[462] = 13'h1066;
        RAM[463] = 13'h1064;
        RAM[464] = 13'h1062;
        RAM[465] = 13'h1060;
        RAM[466] = 13'h105e;
        RAM[467] = 13'h105c;
        RAM[468] = 13'h1059;
        RAM[469] = 13'h1057;
        RAM[470] = 13'h1055;
        RAM[471] = 13'h1053;
        RAM[472] = 13'h1051;
        RAM[473] = 13'h104f;
        RAM[474] = 13'h104d;
        RAM[475] = 13'h104b;
        RAM[476] = 13'h1048;
        RAM[477] = 13'h1046;
        RAM[478] = 13'h1044;
        RAM[479] = 13'h1042;
        RAM[480] = 13'h1040;
        RAM[481] = 13'h103e;
        RAM[482] = 13'h103c;
        RAM[483] = 13'h103a;
        RAM[484] = 13'h1038;
        RAM[485] = 13'h1036;
        RAM[486] = 13'h1033;
        RAM[487] = 13'h1031;
        RAM[488] = 13'h102f;
        RAM[489] = 13'h102d;
        RAM[490] = 13'h102b;
        RAM[491] = 13'h1029;
        RAM[492] = 13'h1027;
        RAM[493] = 13'h1025;
        RAM[494] = 13'h1023;
        RAM[495] = 13'h1021;
        RAM[496] = 13'h101f;
        RAM[497] = 13'h101d;
        RAM[498] = 13'h101b;
        RAM[499] = 13'h1019;
        RAM[500] = 13'h1017;
        RAM[501] = 13'h1015;
        RAM[502] = 13'h1013;
        RAM[503] = 13'h1011;
        RAM[504] = 13'h100f;
        RAM[505] = 13'h100d;
        RAM[506] = 13'h100b;
        RAM[507] = 13'h1009;
        RAM[508] = 13'h1007;
        RAM[509] = 13'h1005;
        RAM[510] = 13'h1003;
        RAM[511] = 13'h1001;
        RAM[512] = 13'h1ffc;
        RAM[513] = 13'h1ff4;
        RAM[514] = 13'h1fec;
        RAM[515] = 13'h1fe4;
        RAM[516] = 13'h1fdc;
        RAM[517] = 13'h1fd4;
        RAM[518] = 13'h1fcc;
        RAM[519] = 13'h1fc4;
        RAM[520] = 13'h1fbc;
        RAM[521] = 13'h1fb5;
        RAM[522] = 13'h1fad;
        RAM[523] = 13'h1fa5;
        RAM[524] = 13'h1f9d;
        RAM[525] = 13'h1f96;
        RAM[526] = 13'h1f8e;
        RAM[527] = 13'h1f86;
        RAM[528] = 13'h1f7f;
        RAM[529] = 13'h1f77;
        RAM[530] = 13'h1f6f;
        RAM[531] = 13'h1f68;
        RAM[532] = 13'h1f60;
        RAM[533] = 13'h1f59;
        RAM[534] = 13'h1f51;
        RAM[535] = 13'h1f4a;
        RAM[536] = 13'h1f42;
        RAM[537] = 13'h1f3b;
        RAM[538] = 13'h1f33;
        RAM[539] = 13'h1f2c;
        RAM[540] = 13'h1f25;
        RAM[541] = 13'h1f1d;
        RAM[542] = 13'h1f16;
        RAM[543] = 13'h1f0f;
        RAM[544] = 13'h1f07;
        RAM[545] = 13'h1f00;
        RAM[546] = 13'h1ef9;
        RAM[547] = 13'h1ef1;
        RAM[548] = 13'h1eea;
        RAM[549] = 13'h1ee3;
        RAM[550] = 13'h1edc;
        RAM[551] = 13'h1ed5;
        RAM[552] = 13'h1ece;
        RAM[553] = 13'h1ec6;
        RAM[554] = 13'h1ebf;
        RAM[555] = 13'h1eb8;
        RAM[556] = 13'h1eb1;
        RAM[557] = 13'h1eaa;
        RAM[558] = 13'h1ea3;
        RAM[559] = 13'h1e9c;
        RAM[560] = 13'h1e95;
        RAM[561] = 13'h1e8e;
        RAM[562] = 13'h1e87;
        RAM[563] = 13'h1e80;
        RAM[564] = 13'h1e79;
        RAM[565] = 13'h1e72;
        RAM[566] = 13'h1e6b;
        RAM[567] = 13'h1e65;
        RAM[568] = 13'h1e5e;
        RAM[569] = 13'h1e57;
        RAM[570] = 13'h1e50;
        RAM[571] = 13'h1e49;
        RAM[572] = 13'h1e43;
        RAM[573] = 13'h1e3c;
        RAM[574] = 13'h1e35;
        RAM[575] = 13'h1e2e;
        RAM[576] = 13'h1e28;
        RAM[577] = 13'h1e21;
        RAM[578] = 13'h1e1a;
        RAM[579] = 13'h1e14;
        RAM[580] = 13'h1e0d;
        RAM[581] = 13'h1e06;
        RAM[582] = 13'h1e00;
        RAM[583] = 13'h1df9;
        RAM[584] = 13'h1df3;
        RAM[585] = 13'h1dec;
        RAM[586] = 13'h1de6;
        RAM[587] = 13'h1ddf;
        RAM[588] = 13'h1dd9;
        RAM[589] = 13'h1dd2;
        RAM[590] = 13'h1dcc;
        RAM[591] = 13'h1dc5;
        RAM[592] = 13'h1dbf;
        RAM[593] = 13'h1db8;
        RAM[594] = 13'h1db2;
        RAM[595] = 13'h1dab;
        RAM[596] = 13'h1da5;
        RAM[597] = 13'h1d9f;
        RAM[598] = 13'h1d98;
        RAM[599] = 13'h1d92;
        RAM[600] = 13'h1d8c;
        RAM[601] = 13'h1d86;
        RAM[602] = 13'h1d7f;
        RAM[603] = 13'h1d79;
        RAM[604] = 13'h1d73;
        RAM[605] = 13'h1d6c;
        RAM[606] = 13'h1d66;
        RAM[607] = 13'h1d60;
        RAM[608] = 13'h1d5a;
        RAM[609] = 13'h1d54;
        RAM[610] = 13'h1d4e;
        RAM[611] = 13'h1d47;
        RAM[612] = 13'h1d41;
        RAM[613] = 13'h1d3b;
        RAM[614] = 13'h1d35;
        RAM[615] = 13'h1d2f;
        RAM[616] = 13'h1d29;
        RAM[617] = 13'h1d23;
        RAM[618] = 13'h1d1d;
        RAM[619] = 13'h1d17;
        RAM[620] = 13'h1d11;
        RAM[621] = 13'h1d0b;
        RAM[622] = 13'h1d05;
        RAM[623] = 13'h1cff;
        RAM[624] = 13'h1cf9;
        RAM[625] = 13'h1cf3;
        RAM[626] = 13'h1ced;
        RAM[627] = 13'h1ce7;
        RAM[628] = 13'h1ce1;
        RAM[629] = 13'h1cdc;
        RAM[630] = 13'h1cd6;
        RAM[631] = 13'h1cd0;
        RAM[632] = 13'h1cca;
        RAM[633] = 13'h1cc4;
        RAM[634] = 13'h1cbe;
        RAM[635] = 13'h1cb9;
        RAM[636] = 13'h1cb3;
        RAM[637] = 13'h1cad;
        RAM[638] = 13'h1ca7;
        RAM[639] = 13'h1ca2;
        RAM[640] = 13'h1c9c;
        RAM[641] = 13'h1c96;
        RAM[642] = 13'h1c90;
        RAM[643] = 13'h1c8b;
        RAM[644] = 13'h1c85;
        RAM[645] = 13'h1c7f;
        RAM[646] = 13'h1c7a;
        RAM[647] = 13'h1c74;
        RAM[648] = 13'h1c6e;
        RAM[649] = 13'h1c69;
        RAM[650] = 13'h1c63;
        RAM[651] = 13'h1c5e;
        RAM[652] = 13'h1c58;
        RAM[653] = 13'h1c53;
        RAM[654] = 13'h1c4d;
        RAM[655] = 13'h1c48;
        RAM[656] = 13'h1c42;
        RAM[657] = 13'h1c3c;
        RAM[658] = 13'h1c37;
        RAM[659] = 13'h1c32;
        RAM[660] = 13'h1c2c;
        RAM[661] = 13'h1c27;
        RAM[662] = 13'h1c21;
        RAM[663] = 13'h1c1c;
        RAM[664] = 13'h1c16;
        RAM[665] = 13'h1c11;
        RAM[666] = 13'h1c0c;
        RAM[667] = 13'h1c06;
        RAM[668] = 13'h1c01;
        RAM[669] = 13'h1bfb;
        RAM[670] = 13'h1bf6;
        RAM[671] = 13'h1bf1;
        RAM[672] = 13'h1beb;
        RAM[673] = 13'h1be6;
        RAM[674] = 13'h1be1;
        RAM[675] = 13'h1bdc;
        RAM[676] = 13'h1bd6;
        RAM[677] = 13'h1bd1;
        RAM[678] = 13'h1bcc;
        RAM[679] = 13'h1bc6;
        RAM[680] = 13'h1bc1;
        RAM[681] = 13'h1bbc;
        RAM[682] = 13'h1bb7;
        RAM[683] = 13'h1bb2;
        RAM[684] = 13'h1bac;
        RAM[685] = 13'h1ba7;
        RAM[686] = 13'h1ba2;
        RAM[687] = 13'h1b9d;
        RAM[688] = 13'h1b98;
        RAM[689] = 13'h1b93;
        RAM[690] = 13'h1b8e;
        RAM[691] = 13'h1b89;
        RAM[692] = 13'h1b83;
        RAM[693] = 13'h1b7e;
        RAM[694] = 13'h1b79;
        RAM[695] = 13'h1b74;
        RAM[696] = 13'h1b6f;
        RAM[697] = 13'h1b6a;
        RAM[698] = 13'h1b65;
        RAM[699] = 13'h1b60;
        RAM[700] = 13'h1b5b;
        RAM[701] = 13'h1b56;
        RAM[702] = 13'h1b51;
        RAM[703] = 13'h1b4c;
        RAM[704] = 13'h1b47;
        RAM[705] = 13'h1b42;
        RAM[706] = 13'h1b3d;
        RAM[707] = 13'h1b38;
        RAM[708] = 13'h1b33;
        RAM[709] = 13'h1b2f;
        RAM[710] = 13'h1b2a;
        RAM[711] = 13'h1b25;
        RAM[712] = 13'h1b20;
        RAM[713] = 13'h1b1b;
        RAM[714] = 13'h1b16;
        RAM[715] = 13'h1b11;
        RAM[716] = 13'h1b0c;
        RAM[717] = 13'h1b08;
        RAM[718] = 13'h1b03;
        RAM[719] = 13'h1afe;
        RAM[720] = 13'h1af9;
        RAM[721] = 13'h1af4;
        RAM[722] = 13'h1af0;
        RAM[723] = 13'h1aeb;
        RAM[724] = 13'h1ae6;
        RAM[725] = 13'h1ae1;
        RAM[726] = 13'h1add;
        RAM[727] = 13'h1ad8;
        RAM[728] = 13'h1ad3;
        RAM[729] = 13'h1ace;
        RAM[730] = 13'h1aca;
        RAM[731] = 13'h1ac5;
        RAM[732] = 13'h1ac0;
        RAM[733] = 13'h1abc;
        RAM[734] = 13'h1ab7;
        RAM[735] = 13'h1ab2;
        RAM[736] = 13'h1aae;
        RAM[737] = 13'h1aa9;
        RAM[738] = 13'h1aa5;
        RAM[739] = 13'h1aa0;
        RAM[740] = 13'h1a9b;
        RAM[741] = 13'h1a97;
        RAM[742] = 13'h1a92;
        RAM[743] = 13'h1a8e;
        RAM[744] = 13'h1a89;
        RAM[745] = 13'h1a84;
        RAM[746] = 13'h1a80;
        RAM[747] = 13'h1a7b;
        RAM[748] = 13'h1a77;
        RAM[749] = 13'h1a72;
        RAM[750] = 13'h1a6e;
        RAM[751] = 13'h1a69;
        RAM[752] = 13'h1a65;
        RAM[753] = 13'h1a60;
        RAM[754] = 13'h1a5c;
        RAM[755] = 13'h1a57;
        RAM[756] = 13'h1a53;
        RAM[757] = 13'h1a4e;
        RAM[758] = 13'h1a4a;
        RAM[759] = 13'h1a46;
        RAM[760] = 13'h1a41;
        RAM[761] = 13'h1a3d;
        RAM[762] = 13'h1a38;
        RAM[763] = 13'h1a34;
        RAM[764] = 13'h1a30;
        RAM[765] = 13'h1a2b;
        RAM[766] = 13'h1a27;
        RAM[767] = 13'h1a22;
        RAM[768] = 13'h1a1e;
        RAM[769] = 13'h1a1a;
        RAM[770] = 13'h1a15;
        RAM[771] = 13'h1a11;
        RAM[772] = 13'h1a0d;
        RAM[773] = 13'h1a08;
        RAM[774] = 13'h1a04;
        RAM[775] = 13'h1a00;
        RAM[776] = 13'h19fc;
        RAM[777] = 13'h19f7;
        RAM[778] = 13'h19f3;
        RAM[779] = 13'h19ef;
        RAM[780] = 13'h19ea;
        RAM[781] = 13'h19e6;
        RAM[782] = 13'h19e2;
        RAM[783] = 13'h19de;
        RAM[784] = 13'h19da;
        RAM[785] = 13'h19d5;
        RAM[786] = 13'h19d1;
        RAM[787] = 13'h19cd;
        RAM[788] = 13'h19c9;
        RAM[789] = 13'h19c5;
        RAM[790] = 13'h19c0;
        RAM[791] = 13'h19bc;
        RAM[792] = 13'h19b8;
        RAM[793] = 13'h19b4;
        RAM[794] = 13'h19b0;
        RAM[795] = 13'h19ac;
        RAM[796] = 13'h19a7;
        RAM[797] = 13'h19a3;
        RAM[798] = 13'h199f;
        RAM[799] = 13'h199b;
        RAM[800] = 13'h1997;
        RAM[801] = 13'h1993;
        RAM[802] = 13'h198f;
        RAM[803] = 13'h198b;
        RAM[804] = 13'h1987;
        RAM[805] = 13'h1983;
        RAM[806] = 13'h197f;
        RAM[807] = 13'h197b;
        RAM[808] = 13'h1977;
        RAM[809] = 13'h1973;
        RAM[810] = 13'h196f;
        RAM[811] = 13'h196a;
        RAM[812] = 13'h1966;
        RAM[813] = 13'h1962;
        RAM[814] = 13'h195f;
        RAM[815] = 13'h195b;
        RAM[816] = 13'h1957;
        RAM[817] = 13'h1953;
        RAM[818] = 13'h194f;
        RAM[819] = 13'h194b;
        RAM[820] = 13'h1947;
        RAM[821] = 13'h1943;
        RAM[822] = 13'h193f;
        RAM[823] = 13'h193b;
        RAM[824] = 13'h1937;
        RAM[825] = 13'h1933;
        RAM[826] = 13'h192f;
        RAM[827] = 13'h192b;
        RAM[828] = 13'h1927;
        RAM[829] = 13'h1924;
        RAM[830] = 13'h1920;
        RAM[831] = 13'h191c;
        RAM[832] = 13'h1918;
        RAM[833] = 13'h1914;
        RAM[834] = 13'h1910;
        RAM[835] = 13'h190c;
        RAM[836] = 13'h1909;
        RAM[837] = 13'h1905;
        RAM[838] = 13'h1901;
        RAM[839] = 13'h18fd;
        RAM[840] = 13'h18f9;
        RAM[841] = 13'h18f5;
        RAM[842] = 13'h18f2;
        RAM[843] = 13'h18ee;
        RAM[844] = 13'h18ea;
        RAM[845] = 13'h18e6;
        RAM[846] = 13'h18e3;
        RAM[847] = 13'h18df;
        RAM[848] = 13'h18db;
        RAM[849] = 13'h18d7;
        RAM[850] = 13'h18d4;
        RAM[851] = 13'h18d0;
        RAM[852] = 13'h18cc;
        RAM[853] = 13'h18c8;
        RAM[854] = 13'h18c5;
        RAM[855] = 13'h18c1;
        RAM[856] = 13'h18bd;
        RAM[857] = 13'h18ba;
        RAM[858] = 13'h18b6;
        RAM[859] = 13'h18b2;
        RAM[860] = 13'h18af;
        RAM[861] = 13'h18ab;
        RAM[862] = 13'h18a7;
        RAM[863] = 13'h18a4;
        RAM[864] = 13'h18a0;
        RAM[865] = 13'h189c;
        RAM[866] = 13'h1899;
        RAM[867] = 13'h1895;
        RAM[868] = 13'h1891;
        RAM[869] = 13'h188e;
        RAM[870] = 13'h188a;
        RAM[871] = 13'h1887;
        RAM[872] = 13'h1883;
        RAM[873] = 13'h187f;
        RAM[874] = 13'h187c;
        RAM[875] = 13'h1878;
        RAM[876] = 13'h1875;
        RAM[877] = 13'h1871;
        RAM[878] = 13'h186d;
        RAM[879] = 13'h186a;
        RAM[880] = 13'h1866;
        RAM[881] = 13'h1863;
        RAM[882] = 13'h185f;
        RAM[883] = 13'h185c;
        RAM[884] = 13'h1858;
        RAM[885] = 13'h1855;
        RAM[886] = 13'h1851;
        RAM[887] = 13'h184e;
        RAM[888] = 13'h184a;
        RAM[889] = 13'h1847;
        RAM[890] = 13'h1843;
        RAM[891] = 13'h1840;
        RAM[892] = 13'h183c;
        RAM[893] = 13'h1839;
        RAM[894] = 13'h1835;
        RAM[895] = 13'h1832;
        RAM[896] = 13'h182e;
        RAM[897] = 13'h182b;
        RAM[898] = 13'h1827;
        RAM[899] = 13'h1824;
        RAM[900] = 13'h1821;
        RAM[901] = 13'h181d;
        RAM[902] = 13'h181a;
        RAM[903] = 13'h1816;
        RAM[904] = 13'h1813;
        RAM[905] = 13'h1810;
        RAM[906] = 13'h180c;
        RAM[907] = 13'h1809;
        RAM[908] = 13'h1805;
        RAM[909] = 13'h1802;
        RAM[910] = 13'h17ff;
        RAM[911] = 13'h17fb;
        RAM[912] = 13'h17f8;
        RAM[913] = 13'h17f4;
        RAM[914] = 13'h17f1;
        RAM[915] = 13'h17ee;
        RAM[916] = 13'h17ea;
        RAM[917] = 13'h17e7;
        RAM[918] = 13'h17e4;
        RAM[919] = 13'h17e0;
        RAM[920] = 13'h17dd;
        RAM[921] = 13'h17da;
        RAM[922] = 13'h17d6;
        RAM[923] = 13'h17d3;
        RAM[924] = 13'h17d0;
        RAM[925] = 13'h17cd;
        RAM[926] = 13'h17c9;
        RAM[927] = 13'h17c6;
        RAM[928] = 13'h17c3;
        RAM[929] = 13'h17bf;
        RAM[930] = 13'h17bc;
        RAM[931] = 13'h17b9;
        RAM[932] = 13'h17b6;
        RAM[933] = 13'h17b2;
        RAM[934] = 13'h17af;
        RAM[935] = 13'h17ac;
        RAM[936] = 13'h17a9;
        RAM[937] = 13'h17a5;
        RAM[938] = 13'h17a2;
        RAM[939] = 13'h179f;
        RAM[940] = 13'h179c;
        RAM[941] = 13'h1799;
        RAM[942] = 13'h1795;
        RAM[943] = 13'h1792;
        RAM[944] = 13'h178f;
        RAM[945] = 13'h178c;
        RAM[946] = 13'h1789;
        RAM[947] = 13'h1785;
        RAM[948] = 13'h1782;
        RAM[949] = 13'h177f;
        RAM[950] = 13'h177c;
        RAM[951] = 13'h1779;
        RAM[952] = 13'h1776;
        RAM[953] = 13'h1772;
        RAM[954] = 13'h176f;
        RAM[955] = 13'h176c;
        RAM[956] = 13'h1769;
        RAM[957] = 13'h1766;
        RAM[958] = 13'h1763;
        RAM[959] = 13'h1760;
        RAM[960] = 13'h175d;
        RAM[961] = 13'h1759;
        RAM[962] = 13'h1756;
        RAM[963] = 13'h1753;
        RAM[964] = 13'h1750;
        RAM[965] = 13'h174d;
        RAM[966] = 13'h174a;
        RAM[967] = 13'h1747;
        RAM[968] = 13'h1744;
        RAM[969] = 13'h1741;
        RAM[970] = 13'h173e;
        RAM[971] = 13'h173b;
        RAM[972] = 13'h1738;
        RAM[973] = 13'h1734;
        RAM[974] = 13'h1731;
        RAM[975] = 13'h172e;
        RAM[976] = 13'h172b;
        RAM[977] = 13'h1728;
        RAM[978] = 13'h1725;
        RAM[979] = 13'h1722;
        RAM[980] = 13'h171f;
        RAM[981] = 13'h171c;
        RAM[982] = 13'h1719;
        RAM[983] = 13'h1716;
        RAM[984] = 13'h1713;
        RAM[985] = 13'h1710;
        RAM[986] = 13'h170d;
        RAM[987] = 13'h170a;
        RAM[988] = 13'h1707;
        RAM[989] = 13'h1704;
        RAM[990] = 13'h1701;
        RAM[991] = 13'h16fe;
        RAM[992] = 13'h16fb;
        RAM[993] = 13'h16f8;
        RAM[994] = 13'h16f5;
        RAM[995] = 13'h16f2;
        RAM[996] = 13'h16f0;
        RAM[997] = 13'h16ed;
        RAM[998] = 13'h16ea;
        RAM[999] = 13'h16e7;
        RAM[1000] = 13'h16e4;
        RAM[1001] = 13'h16e1;
        RAM[1002] = 13'h16de;
        RAM[1003] = 13'h16db;
        RAM[1004] = 13'h16d8;
        RAM[1005] = 13'h16d5;
        RAM[1006] = 13'h16d2;
        RAM[1007] = 13'h16cf;
        RAM[1008] = 13'h16cc;
        RAM[1009] = 13'h16ca;
        RAM[1010] = 13'h16c7;
        RAM[1011] = 13'h16c4;
        RAM[1012] = 13'h16c1;
        RAM[1013] = 13'h16be;
        RAM[1014] = 13'h16bb;
        RAM[1015] = 13'h16b8;
        RAM[1016] = 13'h16b5;
        RAM[1017] = 13'h16b3;
        RAM[1018] = 13'h16b0;
        RAM[1019] = 13'h16ad;
        RAM[1020] = 13'h16aa;
        RAM[1021] = 13'h16a7;
        RAM[1022] = 13'h16a4;
        RAM[1023] = 13'h16a2;
    end
endmodule
`default_nettype wire
