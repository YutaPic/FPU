`default_nettype none
`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Yuta Fukushima
// 
// Create Date: 2020/10/30
// Design Name: finv_table
// Module Name: finv_const_table, finv_grad_table
// Project Name: C&P
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
//////////////////////////////////////////////////////////////////////////////////
// finv_const_table : ニュートン法線形近似の定数項(23bit)
// finv_grad_table : 勾配(13bit)
// それぞれblockRAM を１ずつ使用
module finv_const_table (
    input wire clk, 
    input wire [9:0] addr,
    output reg [22:0] con);

reg [22:0] RAM [1023:0];
always @(posedge clk)
    con <= RAM[addr];
initial begin
    RAM[0] = 23'h7ffffd;
    RAM[1] = 23'h7fc00d;
    RAM[2] = 23'h7f803d;
    RAM[3] = 23'h7f408d;
    RAM[4] = 23'h7f00fc;
    RAM[5] = 23'h7ec18b;
    RAM[6] = 23'h7e823a;
    RAM[7] = 23'h7e4308;
    RAM[8] = 23'h7e03f5;
    RAM[9] = 23'h7dc502;
    RAM[10] = 23'h7d862e;
    RAM[11] = 23'h7d4778;
    RAM[12] = 23'h7d08e2;
    RAM[13] = 23'h7cca6b;
    RAM[14] = 23'h7c8c13;
    RAM[15] = 23'h7c4dd9;
    RAM[16] = 23'h7c0fbe;
    RAM[17] = 23'h7bd1c1;
    RAM[18] = 23'h7b93e3;
    RAM[19] = 23'h7b5624;
    RAM[20] = 23'h7b1882;
    RAM[21] = 23'h7adaff;
    RAM[22] = 23'h7a9d9a;
    RAM[23] = 23'h7a6053;
    RAM[24] = 23'h7a232a;
    RAM[25] = 23'h79e61f;
    RAM[26] = 23'h79a931;
    RAM[27] = 23'h796c61;
    RAM[28] = 23'h792faf;
    RAM[29] = 23'h78f31a;
    RAM[30] = 23'h78b6a3;
    RAM[31] = 23'h787a49;
    RAM[32] = 23'h783e0d;
    RAM[33] = 23'h7801ed;
    RAM[34] = 23'h77c5eb;
    RAM[35] = 23'h778a05;
    RAM[36] = 23'h774e3d;
    RAM[37] = 23'h771291;
    RAM[38] = 23'h76d702;
    RAM[39] = 23'h769b90;
    RAM[40] = 23'h76603b;
    RAM[41] = 23'h762502;
    RAM[42] = 23'h75e9e5;
    RAM[43] = 23'h75aee5;
    RAM[44] = 23'h757401;
    RAM[45] = 23'h753939;
    RAM[46] = 23'h74fe8e;
    RAM[47] = 23'h74c3fe;
    RAM[48] = 23'h74898a;
    RAM[49] = 23'h744f33;
    RAM[50] = 23'h7414f7;
    RAM[51] = 23'h73dad7;
    RAM[52] = 23'h73a0d2;
    RAM[53] = 23'h7366e9;
    RAM[54] = 23'h732d1c;
    RAM[55] = 23'h72f36a;
    RAM[56] = 23'h72b9d3;
    RAM[57] = 23'h728058;
    RAM[58] = 23'h7246f8;
    RAM[59] = 23'h720db3;
    RAM[60] = 23'h71d489;
    RAM[61] = 23'h719b7a;
    RAM[62] = 23'h716286;
    RAM[63] = 23'h7129ad;
    RAM[64] = 23'h70f0ee;
    RAM[65] = 23'h70b84a;
    RAM[66] = 23'h707fc1;
    RAM[67] = 23'h704752;
    RAM[68] = 23'h700efe;
    RAM[69] = 23'h6fd6c4;
    RAM[70] = 23'h6f9ea5;
    RAM[71] = 23'h6f669f;
    RAM[72] = 23'h6f2eb4;
    RAM[73] = 23'h6ef6e3;
    RAM[74] = 23'h6ebf2c;
    RAM[75] = 23'h6e878f;
    RAM[76] = 23'h6e500c;
    RAM[77] = 23'h6e18a3;
    RAM[78] = 23'h6de153;
    RAM[79] = 23'h6daa1d;
    RAM[80] = 23'h6d7301;
    RAM[81] = 23'h6d3bfe;
    RAM[82] = 23'h6d0515;
    RAM[83] = 23'h6cce45;
    RAM[84] = 23'h6c978e;
    RAM[85] = 23'h6c60f1;
    RAM[86] = 23'h6c2a6d;
    RAM[87] = 23'h6bf402;
    RAM[88] = 23'h6bbdb0;
    RAM[89] = 23'h6b8777;
    RAM[90] = 23'h6b5157;
    RAM[91] = 23'h6b1b50;
    RAM[92] = 23'h6ae561;
    RAM[93] = 23'h6aaf8c;
    RAM[94] = 23'h6a79cf;
    RAM[95] = 23'h6a442a;
    RAM[96] = 23'h6a0e9e;
    RAM[97] = 23'h69d92b;
    RAM[98] = 23'h69a3d0;
    RAM[99] = 23'h696e8d;
    RAM[100] = 23'h693963;
    RAM[101] = 23'h690450;
    RAM[102] = 23'h68cf56;
    RAM[103] = 23'h689a74;
    RAM[104] = 23'h6865aa;
    RAM[105] = 23'h6830f8;
    RAM[106] = 23'h67fc5e;
    RAM[107] = 23'h67c7db;
    RAM[108] = 23'h679370;
    RAM[109] = 23'h675f1d;
    RAM[110] = 23'h672ae2;
    RAM[111] = 23'h66f6be;
    RAM[112] = 23'h66c2b2;
    RAM[113] = 23'h668ebd;
    RAM[114] = 23'h665adf;
    RAM[115] = 23'h662719;
    RAM[116] = 23'h65f36a;
    RAM[117] = 23'h65bfd3;
    RAM[118] = 23'h658c52;
    RAM[119] = 23'h6558e8;
    RAM[120] = 23'h652596;
    RAM[121] = 23'h64f25a;
    RAM[122] = 23'h64bf35;
    RAM[123] = 23'h648c28;
    RAM[124] = 23'h645931;
    RAM[125] = 23'h642650;
    RAM[126] = 23'h63f386;
    RAM[127] = 23'h63c0d3;
    RAM[128] = 23'h638e37;
    RAM[129] = 23'h635bb0;
    RAM[130] = 23'h632941;
    RAM[131] = 23'h62f6e7;
    RAM[132] = 23'h62c4a4;
    RAM[133] = 23'h629277;
    RAM[134] = 23'h626061;
    RAM[135] = 23'h622e60;
    RAM[136] = 23'h61fc76;
    RAM[137] = 23'h61caa1;
    RAM[138] = 23'h6198e3;
    RAM[139] = 23'h61673a;
    RAM[140] = 23'h6135a8;
    RAM[141] = 23'h61042b;
    RAM[142] = 23'h60d2c3;
    RAM[143] = 23'h60a172;
    RAM[144] = 23'h607036;
    RAM[145] = 23'h603f10;
    RAM[146] = 23'h600dff;
    RAM[147] = 23'h5fdd03;
    RAM[148] = 23'h5fac1d;
    RAM[149] = 23'h5f7b4d;
    RAM[150] = 23'h5f4a91;
    RAM[151] = 23'h5f19eb;
    RAM[152] = 23'h5ee95a;
    RAM[153] = 23'h5eb8de;
    RAM[154] = 23'h5e8878;
    RAM[155] = 23'h5e5826;
    RAM[156] = 23'h5e27e9;
    RAM[157] = 23'h5df7c1;
    RAM[158] = 23'h5dc7ae;
    RAM[159] = 23'h5d97b0;
    RAM[160] = 23'h5d67c7;
    RAM[161] = 23'h5d37f2;
    RAM[162] = 23'h5d0832;
    RAM[163] = 23'h5cd886;
    RAM[164] = 23'h5ca8ef;
    RAM[165] = 23'h5c796d;
    RAM[166] = 23'h5c49ff;
    RAM[167] = 23'h5c1aa5;
    RAM[168] = 23'h5beb60;
    RAM[169] = 23'h5bbc2f;
    RAM[170] = 23'h5b8d12;
    RAM[171] = 23'h5b5e0a;
    RAM[172] = 23'h5b2f15;
    RAM[173] = 23'h5b0035;
    RAM[174] = 23'h5ad168;
    RAM[175] = 23'h5aa2b0;
    RAM[176] = 23'h5a740c;
    RAM[177] = 23'h5a457b;
    RAM[178] = 23'h5a16fe;
    RAM[179] = 23'h59e896;
    RAM[180] = 23'h59ba40;
    RAM[181] = 23'h598bff;
    RAM[182] = 23'h595dd1;
    RAM[183] = 23'h592fb7;
    RAM[184] = 23'h5901b0;
    RAM[185] = 23'h58d3bd;
    RAM[186] = 23'h58a5dd;
    RAM[187] = 23'h587811;
    RAM[188] = 23'h584a58;
    RAM[189] = 23'h581cb2;
    RAM[190] = 23'h57ef1f;
    RAM[191] = 23'h57c1a0;
    RAM[192] = 23'h579434;
    RAM[193] = 23'h5766db;
    RAM[194] = 23'h573995;
    RAM[195] = 23'h570c62;
    RAM[196] = 23'h56df42;
    RAM[197] = 23'h56b235;
    RAM[198] = 23'h56853b;
    RAM[199] = 23'h565854;
    RAM[200] = 23'h562b7f;
    RAM[201] = 23'h55febd;
    RAM[202] = 23'h55d20e;
    RAM[203] = 23'h55a572;
    RAM[204] = 23'h5578e8;
    RAM[205] = 23'h554c70;
    RAM[206] = 23'h55200c;
    RAM[207] = 23'h54f3b9;
    RAM[208] = 23'h54c779;
    RAM[209] = 23'h549b4c;
    RAM[210] = 23'h546f30;
    RAM[211] = 23'h544327;
    RAM[212] = 23'h541731;
    RAM[213] = 23'h53eb4c;
    RAM[214] = 23'h53bf7a;
    RAM[215] = 23'h5393ba;
    RAM[216] = 23'h53680b;
    RAM[217] = 23'h533c6f;
    RAM[218] = 23'h5310e5;
    RAM[219] = 23'h52e56d;
    RAM[220] = 23'h52ba07;
    RAM[221] = 23'h528eb2;
    RAM[222] = 23'h52636f;
    RAM[223] = 23'h52383e;
    RAM[224] = 23'h520d1f;
    RAM[225] = 23'h51e212;
    RAM[226] = 23'h51b716;
    RAM[227] = 23'h518c2b;
    RAM[228] = 23'h516153;
    RAM[229] = 23'h51368b;
    RAM[230] = 23'h510bd5;
    RAM[231] = 23'h50e131;
    RAM[232] = 23'h50b69e;
    RAM[233] = 23'h508c1c;
    RAM[234] = 23'h5061ac;
    RAM[235] = 23'h50374d;
    RAM[236] = 23'h500cff;
    RAM[237] = 23'h4fe2c2;
    RAM[238] = 23'h4fb897;
    RAM[239] = 23'h4f8e7c;
    RAM[240] = 23'h4f6473;
    RAM[241] = 23'h4f3a7b;
    RAM[242] = 23'h4f1093;
    RAM[243] = 23'h4ee6bd;
    RAM[244] = 23'h4ebcf7;
    RAM[245] = 23'h4e9342;
    RAM[246] = 23'h4e699e;
    RAM[247] = 23'h4e400b;
    RAM[248] = 23'h4e1689;
    RAM[249] = 23'h4ded17;
    RAM[250] = 23'h4dc3b6;
    RAM[251] = 23'h4d9a66;
    RAM[252] = 23'h4d7126;
    RAM[253] = 23'h4d47f6;
    RAM[254] = 23'h4d1ed8;
    RAM[255] = 23'h4cf5c9;
    RAM[256] = 23'h4ccccb;
    RAM[257] = 23'h4ca3de;
    RAM[258] = 23'h4c7b00;
    RAM[259] = 23'h4c5234;
    RAM[260] = 23'h4c2977;
    RAM[261] = 23'h4c00ca;
    RAM[262] = 23'h4bd82e;
    RAM[263] = 23'h4bafa2;
    RAM[264] = 23'h4b8726;
    RAM[265] = 23'h4b5eba;
    RAM[266] = 23'h4b365f;
    RAM[267] = 23'h4b0e13;
    RAM[268] = 23'h4ae5d7;
    RAM[269] = 23'h4abdab;
    RAM[270] = 23'h4a958f;
    RAM[271] = 23'h4a6d83;
    RAM[272] = 23'h4a4586;
    RAM[273] = 23'h4a1d9a;
    RAM[274] = 23'h49f5bd;
    RAM[275] = 23'h49cdf0;
    RAM[276] = 23'h49a633;
    RAM[277] = 23'h497e85;
    RAM[278] = 23'h4956e7;
    RAM[279] = 23'h492f58;
    RAM[280] = 23'h4907d9;
    RAM[281] = 23'h48e069;
    RAM[282] = 23'h48b909;
    RAM[283] = 23'h4891b8;
    RAM[284] = 23'h486a77;
    RAM[285] = 23'h484345;
    RAM[286] = 23'h481c23;
    RAM[287] = 23'h47f50f;
    RAM[288] = 23'h47ce0b;
    RAM[289] = 23'h47a716;
    RAM[290] = 23'h478030;
    RAM[291] = 23'h47595a;
    RAM[292] = 23'h473292;
    RAM[293] = 23'h470bda;
    RAM[294] = 23'h46e531;
    RAM[295] = 23'h46be96;
    RAM[296] = 23'h46980b;
    RAM[297] = 23'h46718f;
    RAM[298] = 23'h464b21;
    RAM[299] = 23'h4624c2;
    RAM[300] = 23'h45fe73;
    RAM[301] = 23'h45d832;
    RAM[302] = 23'h45b1ff;
    RAM[303] = 23'h458bdc;
    RAM[304] = 23'h4565c7;
    RAM[305] = 23'h453fc1;
    RAM[306] = 23'h4519ca;
    RAM[307] = 23'h44f3e1;
    RAM[308] = 23'h44ce06;
    RAM[309] = 23'h44a83b;
    RAM[310] = 23'h44827d;
    RAM[311] = 23'h445ccf;
    RAM[312] = 23'h44372e;
    RAM[313] = 23'h44119c;
    RAM[314] = 23'h43ec19;
    RAM[315] = 23'h43c6a4;
    RAM[316] = 23'h43a13d;
    RAM[317] = 23'h437be4;
    RAM[318] = 23'h43569a;
    RAM[319] = 23'h43315d;
    RAM[320] = 23'h430c2f;
    RAM[321] = 23'h42e710;
    RAM[322] = 23'h42c1fe;
    RAM[323] = 23'h429cfa;
    RAM[324] = 23'h427805;
    RAM[325] = 23'h42531d;
    RAM[326] = 23'h422e44;
    RAM[327] = 23'h420978;
    RAM[328] = 23'h41e4bb;
    RAM[329] = 23'h41c00b;
    RAM[330] = 23'h419b69;
    RAM[331] = 23'h4176d5;
    RAM[332] = 23'h41524f;
    RAM[333] = 23'h412dd6;
    RAM[334] = 23'h41096c;
    RAM[335] = 23'h40e50f;
    RAM[336] = 23'h40c0c0;
    RAM[337] = 23'h409c7e;
    RAM[338] = 23'h40784a;
    RAM[339] = 23'h405424;
    RAM[340] = 23'h40300b;
    RAM[341] = 23'h400c00;
    RAM[342] = 23'h3fe802;
    RAM[343] = 23'h3fc412;
    RAM[344] = 23'h3fa02f;
    RAM[345] = 23'h3f7c59;
    RAM[346] = 23'h3f5891;
    RAM[347] = 23'h3f34d7;
    RAM[348] = 23'h3f1129;
    RAM[349] = 23'h3eed89;
    RAM[350] = 23'h3ec9f7;
    RAM[351] = 23'h3ea671;
    RAM[352] = 23'h3e82f9;
    RAM[353] = 23'h3e5f8e;
    RAM[354] = 23'h3e3c30;
    RAM[355] = 23'h3e18df;
    RAM[356] = 23'h3df59b;
    RAM[357] = 23'h3dd265;
    RAM[358] = 23'h3daf3b;
    RAM[359] = 23'h3d8c1f;
    RAM[360] = 23'h3d690f;
    RAM[361] = 23'h3d460d;
    RAM[362] = 23'h3d2317;
    RAM[363] = 23'h3d002e;
    RAM[364] = 23'h3cdd52;
    RAM[365] = 23'h3cba83;
    RAM[366] = 23'h3c97c1;
    RAM[367] = 23'h3c750c;
    RAM[368] = 23'h3c5263;
    RAM[369] = 23'h3c2fc7;
    RAM[370] = 23'h3c0d38;
    RAM[371] = 23'h3beab5;
    RAM[372] = 23'h3bc83f;
    RAM[373] = 23'h3ba5d6;
    RAM[374] = 23'h3b837a;
    RAM[375] = 23'h3b612a;
    RAM[376] = 23'h3b3ee6;
    RAM[377] = 23'h3b1caf;
    RAM[378] = 23'h3afa85;
    RAM[379] = 23'h3ad867;
    RAM[380] = 23'h3ab655;
    RAM[381] = 23'h3a9450;
    RAM[382] = 23'h3a7257;
    RAM[383] = 23'h3a506b;
    RAM[384] = 23'h3a2e8b;
    RAM[385] = 23'h3a0cb7;
    RAM[386] = 23'h39eaef;
    RAM[387] = 23'h39c934;
    RAM[388] = 23'h39a785;
    RAM[389] = 23'h3985e2;
    RAM[390] = 23'h39644c;
    RAM[391] = 23'h3942c1;
    RAM[392] = 23'h392143;
    RAM[393] = 23'h38ffd1;
    RAM[394] = 23'h38de6b;
    RAM[395] = 23'h38bd10;
    RAM[396] = 23'h389bc2;
    RAM[397] = 23'h387a80;
    RAM[398] = 23'h38594a;
    RAM[399] = 23'h383820;
    RAM[400] = 23'h381702;
    RAM[401] = 23'h37f5f0;
    RAM[402] = 23'h37d4e9;
    RAM[403] = 23'h37b3ef;
    RAM[404] = 23'h379300;
    RAM[405] = 23'h37721d;
    RAM[406] = 23'h375146;
    RAM[407] = 23'h37307a;
    RAM[408] = 23'h370fba;
    RAM[409] = 23'h36ef06;
    RAM[410] = 23'h36ce5e;
    RAM[411] = 23'h36adc1;
    RAM[412] = 23'h368d30;
    RAM[413] = 23'h366cab;
    RAM[414] = 23'h364c31;
    RAM[415] = 23'h362bc3;
    RAM[416] = 23'h360b60;
    RAM[417] = 23'h35eb08;
    RAM[418] = 23'h35cabd;
    RAM[419] = 23'h35aa7c;
    RAM[420] = 23'h358a47;
    RAM[421] = 23'h356a1e;
    RAM[422] = 23'h354a00;
    RAM[423] = 23'h3529ed;
    RAM[424] = 23'h3509e6;
    RAM[425] = 23'h34e9ea;
    RAM[426] = 23'h34c9f9;
    RAM[427] = 23'h34aa13;
    RAM[428] = 23'h348a39;
    RAM[429] = 23'h346a6a;
    RAM[430] = 23'h344aa6;
    RAM[431] = 23'h342aed;
    RAM[432] = 23'h340b40;
    RAM[433] = 23'h33eb9d;
    RAM[434] = 23'h33cc06;
    RAM[435] = 23'h33ac7a;
    RAM[436] = 23'h338cf9;
    RAM[437] = 23'h336d83;
    RAM[438] = 23'h334e18;
    RAM[439] = 23'h332eb8;
    RAM[440] = 23'h330f62;
    RAM[441] = 23'h32f018;
    RAM[442] = 23'h32d0d9;
    RAM[443] = 23'h32b1a5;
    RAM[444] = 23'h32927b;
    RAM[445] = 23'h32735d;
    RAM[446] = 23'h325449;
    RAM[447] = 23'h323540;
    RAM[448] = 23'h321642;
    RAM[449] = 23'h31f74f;
    RAM[450] = 23'h31d866;
    RAM[451] = 23'h31b988;
    RAM[452] = 23'h319ab5;
    RAM[453] = 23'h317bec;
    RAM[454] = 23'h315d2f;
    RAM[455] = 23'h313e7b;
    RAM[456] = 23'h311fd3;
    RAM[457] = 23'h310135;
    RAM[458] = 23'h30e2a2;
    RAM[459] = 23'h30c419;
    RAM[460] = 23'h30a59a;
    RAM[461] = 23'h308727;
    RAM[462] = 23'h3068bd;
    RAM[463] = 23'h304a5f;
    RAM[464] = 23'h302c0a;
    RAM[465] = 23'h300dc0;
    RAM[466] = 23'h2fef81;
    RAM[467] = 23'h2fd14c;
    RAM[468] = 23'h2fb321;
    RAM[469] = 23'h2f9500;
    RAM[470] = 23'h2f76ea;
    RAM[471] = 23'h2f58df;
    RAM[472] = 23'h2f3add;
    RAM[473] = 23'h2f1ce6;
    RAM[474] = 23'h2efef9;
    RAM[475] = 23'h2ee116;
    RAM[476] = 23'h2ec33d;
    RAM[477] = 23'h2ea56f;
    RAM[478] = 23'h2e87ab;
    RAM[479] = 23'h2e69f1;
    RAM[480] = 23'h2e4c41;
    RAM[481] = 23'h2e2e9b;
    RAM[482] = 23'h2e10ff;
    RAM[483] = 23'h2df36d;
    RAM[484] = 23'h2dd5e5;
    RAM[485] = 23'h2db868;
    RAM[486] = 23'h2d9af4;
    RAM[487] = 23'h2d7d8a;
    RAM[488] = 23'h2d602b;
    RAM[489] = 23'h2d42d5;
    RAM[490] = 23'h2d2589;
    RAM[491] = 23'h2d0847;
    RAM[492] = 23'h2ceb0f;
    RAM[493] = 23'h2ccde1;
    RAM[494] = 23'h2cb0bc;
    RAM[495] = 23'h2c93a2;
    RAM[496] = 23'h2c7691;
    RAM[497] = 23'h2c598a;
    RAM[498] = 23'h2c3c8d;
    RAM[499] = 23'h2c1f99;
    RAM[500] = 23'h2c02af;
    RAM[501] = 23'h2be5cf;
    RAM[502] = 23'h2bc8f9;
    RAM[503] = 23'h2bac2c;
    RAM[504] = 23'h2b8f69;
    RAM[505] = 23'h2b72b0;
    RAM[506] = 23'h2b5600;
    RAM[507] = 23'h2b395a;
    RAM[508] = 23'h2b1cbd;
    RAM[509] = 23'h2b002a;
    RAM[510] = 23'h2ae3a1;
    RAM[511] = 23'h2ac721;
    RAM[512] = 23'h2aaaaa;
    RAM[513] = 23'h2a8e3d;
    RAM[514] = 23'h2a71d9;
    RAM[515] = 23'h2a557f;
    RAM[516] = 23'h2a392f;
    RAM[517] = 23'h2a1ce7;
    RAM[518] = 23'h2a00a9;
    RAM[519] = 23'h29e475;
    RAM[520] = 23'h29c84a;
    RAM[521] = 23'h29ac28;
    RAM[522] = 23'h29900f;
    RAM[523] = 23'h297400;
    RAM[524] = 23'h2957fa;
    RAM[525] = 23'h293bfd;
    RAM[526] = 23'h29200a;
    RAM[527] = 23'h290420;
    RAM[528] = 23'h28e83f;
    RAM[529] = 23'h28cc67;
    RAM[530] = 23'h28b098;
    RAM[531] = 23'h2894d3;
    RAM[532] = 23'h287916;
    RAM[533] = 23'h285d63;
    RAM[534] = 23'h2841b9;
    RAM[535] = 23'h282618;
    RAM[536] = 23'h280a80;
    RAM[537] = 23'h27eef1;
    RAM[538] = 23'h27d36b;
    RAM[539] = 23'h27b7ee;
    RAM[540] = 23'h279c7a;
    RAM[541] = 23'h278110;
    RAM[542] = 23'h2765ae;
    RAM[543] = 23'h274a55;
    RAM[544] = 23'h272f05;
    RAM[545] = 23'h2713bd;
    RAM[546] = 23'h26f87f;
    RAM[547] = 23'h26dd4a;
    RAM[548] = 23'h26c21d;
    RAM[549] = 23'h26a6fa;
    RAM[550] = 23'h268bdf;
    RAM[551] = 23'h2670cd;
    RAM[552] = 23'h2655c4;
    RAM[553] = 23'h263ac3;
    RAM[554] = 23'h261fcb;
    RAM[555] = 23'h2604dd;
    RAM[556] = 23'h25e9f6;
    RAM[557] = 23'h25cf19;
    RAM[558] = 23'h25b444;
    RAM[559] = 23'h259978;
    RAM[560] = 23'h257eb4;
    RAM[561] = 23'h2563fa;
    RAM[562] = 23'h254947;
    RAM[563] = 23'h252e9e;
    RAM[564] = 23'h2513fd;
    RAM[565] = 23'h24f964;
    RAM[566] = 23'h24ded5;
    RAM[567] = 23'h24c44d;
    RAM[568] = 23'h24a9cf;
    RAM[569] = 23'h248f58;
    RAM[570] = 23'h2474eb;
    RAM[571] = 23'h245a85;
    RAM[572] = 23'h244029;
    RAM[573] = 23'h2425d4;
    RAM[574] = 23'h240b88;
    RAM[575] = 23'h23f145;
    RAM[576] = 23'h23d70a;
    RAM[577] = 23'h23bcd7;
    RAM[578] = 23'h23a2ad;
    RAM[579] = 23'h23888b;
    RAM[580] = 23'h236e71;
    RAM[581] = 23'h235460;
    RAM[582] = 23'h233a57;
    RAM[583] = 23'h232056;
    RAM[584] = 23'h23065e;
    RAM[585] = 23'h22ec6e;
    RAM[586] = 23'h22d286;
    RAM[587] = 23'h22b8a6;
    RAM[588] = 23'h229ecf;
    RAM[589] = 23'h2284ff;
    RAM[590] = 23'h226b38;
    RAM[591] = 23'h225179;
    RAM[592] = 23'h2237c3;
    RAM[593] = 23'h221e14;
    RAM[594] = 23'h22046e;
    RAM[595] = 23'h21eacf;
    RAM[596] = 23'h21d139;
    RAM[597] = 23'h21b7ab;
    RAM[598] = 23'h219e25;
    RAM[599] = 23'h2184a7;
    RAM[600] = 23'h216b31;
    RAM[601] = 23'h2151c3;
    RAM[602] = 23'h21385d;
    RAM[603] = 23'h211eff;
    RAM[604] = 23'h2105a9;
    RAM[605] = 23'h20ec5b;
    RAM[606] = 23'h20d315;
    RAM[607] = 23'h20b9d6;
    RAM[608] = 23'h20a0a0;
    RAM[609] = 23'h208772;
    RAM[610] = 23'h206e4b;
    RAM[611] = 23'h20552d;
    RAM[612] = 23'h203c16;
    RAM[613] = 23'h202307;
    RAM[614] = 23'h200a00;
    RAM[615] = 23'h1ff101;
    RAM[616] = 23'h1fd80a;
    RAM[617] = 23'h1fbf1a;
    RAM[618] = 23'h1fa632;
    RAM[619] = 23'h1f8d52;
    RAM[620] = 23'h1f747a;
    RAM[621] = 23'h1f5ba9;
    RAM[622] = 23'h1f42e0;
    RAM[623] = 23'h1f2a1f;
    RAM[624] = 23'h1f1165;
    RAM[625] = 23'h1ef8b4;
    RAM[626] = 23'h1ee009;
    RAM[627] = 23'h1ec767;
    RAM[628] = 23'h1eaecc;
    RAM[629] = 23'h1e9639;
    RAM[630] = 23'h1e7dad;
    RAM[631] = 23'h1e6529;
    RAM[632] = 23'h1e4cad;
    RAM[633] = 23'h1e3438;
    RAM[634] = 23'h1e1bca;
    RAM[635] = 23'h1e0365;
    RAM[636] = 23'h1deb06;
    RAM[637] = 23'h1dd2b0;
    RAM[638] = 23'h1dba60;
    RAM[639] = 23'h1da219;
    RAM[640] = 23'h1d89d8;
    RAM[641] = 23'h1d719f;
    RAM[642] = 23'h1d596e;
    RAM[643] = 23'h1d4144;
    RAM[644] = 23'h1d2921;
    RAM[645] = 23'h1d1106;
    RAM[646] = 23'h1cf8f2;
    RAM[647] = 23'h1ce0e6;
    RAM[648] = 23'h1cc8e1;
    RAM[649] = 23'h1cb0e3;
    RAM[650] = 23'h1c98ed;
    RAM[651] = 23'h1c80fe;
    RAM[652] = 23'h1c6916;
    RAM[653] = 23'h1c5136;
    RAM[654] = 23'h1c395d;
    RAM[655] = 23'h1c218b;
    RAM[656] = 23'h1c09c0;
    RAM[657] = 23'h1bf1fd;
    RAM[658] = 23'h1bda41;
    RAM[659] = 23'h1bc28c;
    RAM[660] = 23'h1baade;
    RAM[661] = 23'h1b9338;
    RAM[662] = 23'h1b7b98;
    RAM[663] = 23'h1b6400;
    RAM[664] = 23'h1b4c6f;
    RAM[665] = 23'h1b34e5;
    RAM[666] = 23'h1b1d63;
    RAM[667] = 23'h1b05e7;
    RAM[668] = 23'h1aee73;
    RAM[669] = 23'h1ad705;
    RAM[670] = 23'h1abf9f;
    RAM[671] = 23'h1aa840;
    RAM[672] = 23'h1a90e7;
    RAM[673] = 23'h1a7996;
    RAM[674] = 23'h1a624c;
    RAM[675] = 23'h1a4b09;
    RAM[676] = 23'h1a33cd;
    RAM[677] = 23'h1a1c98;
    RAM[678] = 23'h1a056a;
    RAM[679] = 23'h19ee43;
    RAM[680] = 23'h19d722;
    RAM[681] = 23'h19c009;
    RAM[682] = 23'h19a8f7;
    RAM[683] = 23'h1991ec;
    RAM[684] = 23'h197ae7;
    RAM[685] = 23'h1963e9;
    RAM[686] = 23'h194cf3;
    RAM[687] = 23'h193603;
    RAM[688] = 23'h191f1a;
    RAM[689] = 23'h190838;
    RAM[690] = 23'h18f15d;
    RAM[691] = 23'h18da88;
    RAM[692] = 23'h18c3ba;
    RAM[693] = 23'h18acf4;
    RAM[694] = 23'h189634;
    RAM[695] = 23'h187f7a;
    RAM[696] = 23'h1868c8;
    RAM[697] = 23'h18521c;
    RAM[698] = 23'h183b77;
    RAM[699] = 23'h1824d9;
    RAM[700] = 23'h180e41;
    RAM[701] = 23'h17f7b0;
    RAM[702] = 23'h17e126;
    RAM[703] = 23'h17caa2;
    RAM[704] = 23'h17b426;
    RAM[705] = 23'h179daf;
    RAM[706] = 23'h178740;
    RAM[707] = 23'h1770d7;
    RAM[708] = 23'h175a75;
    RAM[709] = 23'h174419;
    RAM[710] = 23'h172dc4;
    RAM[711] = 23'h171776;
    RAM[712] = 23'h17012e;
    RAM[713] = 23'h16eaec;
    RAM[714] = 23'h16d4b2;
    RAM[715] = 23'h16be7d;
    RAM[716] = 23'h16a850;
    RAM[717] = 23'h169229;
    RAM[718] = 23'h167c08;
    RAM[719] = 23'h1665ee;
    RAM[720] = 23'h164fda;
    RAM[721] = 23'h1639cd;
    RAM[722] = 23'h1623c6;
    RAM[723] = 23'h160dc6;
    RAM[724] = 23'h15f7cc;
    RAM[725] = 23'h15e1d9;
    RAM[726] = 23'h15cbec;
    RAM[727] = 23'h15b605;
    RAM[728] = 23'h15a025;
    RAM[729] = 23'h158a4b;
    RAM[730] = 23'h157478;
    RAM[731] = 23'h155eab;
    RAM[732] = 23'h1548e4;
    RAM[733] = 23'h153324;
    RAM[734] = 23'h151d6a;
    RAM[735] = 23'h1507b6;
    RAM[736] = 23'h14f209;
    RAM[737] = 23'h14dc62;
    RAM[738] = 23'h14c6c1;
    RAM[739] = 23'h14b127;
    RAM[740] = 23'h149b93;
    RAM[741] = 23'h148605;
    RAM[742] = 23'h14707d;
    RAM[743] = 23'h145afc;
    RAM[744] = 23'h144580;
    RAM[745] = 23'h14300b;
    RAM[746] = 23'h141a9d;
    RAM[747] = 23'h140534;
    RAM[748] = 23'h13efd1;
    RAM[749] = 23'h13da75;
    RAM[750] = 23'h13c51f;
    RAM[751] = 23'h13afcf;
    RAM[752] = 23'h139a85;
    RAM[753] = 23'h138542;
    RAM[754] = 23'h137004;
    RAM[755] = 23'h135acd;
    RAM[756] = 23'h13459c;
    RAM[757] = 23'h133070;
    RAM[758] = 23'h131b4b;
    RAM[759] = 23'h13062c;
    RAM[760] = 23'h12f113;
    RAM[761] = 23'h12dc00;
    RAM[762] = 23'h12c6f3;
    RAM[763] = 23'h12b1ed;
    RAM[764] = 23'h129cec;
    RAM[765] = 23'h1287f1;
    RAM[766] = 23'h1272fc;
    RAM[767] = 23'h125e0d;
    RAM[768] = 23'h124924;
    RAM[769] = 23'h123441;
    RAM[770] = 23'h121f65;
    RAM[771] = 23'h120a8e;
    RAM[772] = 23'h11f5bc;
    RAM[773] = 23'h11e0f1;
    RAM[774] = 23'h11cc2c;
    RAM[775] = 23'h11b76d;
    RAM[776] = 23'h11a2b4;
    RAM[777] = 23'h118e00;
    RAM[778] = 23'h117952;
    RAM[779] = 23'h1164ab;
    RAM[780] = 23'h115009;
    RAM[781] = 23'h113b6d;
    RAM[782] = 23'h1126d7;
    RAM[783] = 23'h111246;
    RAM[784] = 23'h10fdbc;
    RAM[785] = 23'h10e937;
    RAM[786] = 23'h10d4b8;
    RAM[787] = 23'h10c03f;
    RAM[788] = 23'h10abcc;
    RAM[789] = 23'h10975e;
    RAM[790] = 23'h1082f6;
    RAM[791] = 23'h106e94;
    RAM[792] = 23'h105a38;
    RAM[793] = 23'h1045e2;
    RAM[794] = 23'h103191;
    RAM[795] = 23'h101d46;
    RAM[796] = 23'h100900;
    RAM[797] = 23'hff4c1;
    RAM[798] = 23'hfe087;
    RAM[799] = 23'hfcc52;
    RAM[800] = 23'hfb824;
    RAM[801] = 23'hfa3fb;
    RAM[802] = 23'hf8fd7;
    RAM[803] = 23'hf7bba;
    RAM[804] = 23'hf67a2;
    RAM[805] = 23'hf538f;
    RAM[806] = 23'hf3f82;
    RAM[807] = 23'hf2b7b;
    RAM[808] = 23'hf177a;
    RAM[809] = 23'hf037e;
    RAM[810] = 23'heef87;
    RAM[811] = 23'hedb96;
    RAM[812] = 23'hec7ab;
    RAM[813] = 23'heb3c5;
    RAM[814] = 23'he9fe5;
    RAM[815] = 23'he8c0a;
    RAM[816] = 23'he7835;
    RAM[817] = 23'he6466;
    RAM[818] = 23'he509b;
    RAM[819] = 23'he3cd7;
    RAM[820] = 23'he2918;
    RAM[821] = 23'he155e;
    RAM[822] = 23'he01aa;
    RAM[823] = 23'hdedfb;
    RAM[824] = 23'hdda52;
    RAM[825] = 23'hdc6ae;
    RAM[826] = 23'hdb310;
    RAM[827] = 23'hd9f77;
    RAM[828] = 23'hd8be3;
    RAM[829] = 23'hd7855;
    RAM[830] = 23'hd64cc;
    RAM[831] = 23'hd5149;
    RAM[832] = 23'hd3dcb;
    RAM[833] = 23'hd2a52;
    RAM[834] = 23'hd16df;
    RAM[835] = 23'hd0371;
    RAM[836] = 23'hcf009;
    RAM[837] = 23'hcdca5;
    RAM[838] = 23'hcc948;
    RAM[839] = 23'hcb5ef;
    RAM[840] = 23'hca29c;
    RAM[841] = 23'hc8f4e;
    RAM[842] = 23'hc7c05;
    RAM[843] = 23'hc68c2;
    RAM[844] = 23'hc5584;
    RAM[845] = 23'hc424b;
    RAM[846] = 23'hc2f18;
    RAM[847] = 23'hc1be9;
    RAM[848] = 23'hc08c0;
    RAM[849] = 23'hbf59d;
    RAM[850] = 23'hbe27e;
    RAM[851] = 23'hbcf65;
    RAM[852] = 23'hbbc51;
    RAM[853] = 23'hba942;
    RAM[854] = 23'hb9638;
    RAM[855] = 23'hb8333;
    RAM[856] = 23'hb7034;
    RAM[857] = 23'hb5d3a;
    RAM[858] = 23'hb4a45;
    RAM[859] = 23'hb3755;
    RAM[860] = 23'hb246a;
    RAM[861] = 23'hb1185;
    RAM[862] = 23'hafea4;
    RAM[863] = 23'haebc9;
    RAM[864] = 23'had8f3;
    RAM[865] = 23'hac622;
    RAM[866] = 23'hab356;
    RAM[867] = 23'haa08f;
    RAM[868] = 23'ha8dcd;
    RAM[869] = 23'ha7b10;
    RAM[870] = 23'ha6859;
    RAM[871] = 23'ha55a6;
    RAM[872] = 23'ha42f8;
    RAM[873] = 23'ha3050;
    RAM[874] = 23'ha1dac;
    RAM[875] = 23'ha0b0e;
    RAM[876] = 23'h9f874;
    RAM[877] = 23'h9e5e0;
    RAM[878] = 23'h9d350;
    RAM[879] = 23'h9c0c6;
    RAM[880] = 23'h9ae40;
    RAM[881] = 23'h99bc0;
    RAM[882] = 23'h98944;
    RAM[883] = 23'h976ce;
    RAM[884] = 23'h9645c;
    RAM[885] = 23'h951f0;
    RAM[886] = 23'h93f88;
    RAM[887] = 23'h92d25;
    RAM[888] = 23'h91ac7;
    RAM[889] = 23'h9086e;
    RAM[890] = 23'h8f61a;
    RAM[891] = 23'h8e3cb;
    RAM[892] = 23'h8d181;
    RAM[893] = 23'h8bf3b;
    RAM[894] = 23'h8acfb;
    RAM[895] = 23'h89abf;
    RAM[896] = 23'h88888;
    RAM[897] = 23'h87657;
    RAM[898] = 23'h86429;
    RAM[899] = 23'h85201;
    RAM[900] = 23'h83fde;
    RAM[901] = 23'h82dbf;
    RAM[902] = 23'h81ba6;
    RAM[903] = 23'h80991;
    RAM[904] = 23'h7f780;
    RAM[905] = 23'h7e575;
    RAM[906] = 23'h7d36f;
    RAM[907] = 23'h7c16d;
    RAM[908] = 23'h7af70;
    RAM[909] = 23'h79d77;
    RAM[910] = 23'h78b84;
    RAM[911] = 23'h77995;
    RAM[912] = 23'h767ab;
    RAM[913] = 23'h755c6;
    RAM[914] = 23'h743e5;
    RAM[915] = 23'h7320a;
    RAM[916] = 23'h72033;
    RAM[917] = 23'h70e60;
    RAM[918] = 23'h6fc93;
    RAM[919] = 23'h6eaca;
    RAM[920] = 23'h6d905;
    RAM[921] = 23'h6c746;
    RAM[922] = 23'h6b58b;
    RAM[923] = 23'h6a3d4;
    RAM[924] = 23'h69223;
    RAM[925] = 23'h68076;
    RAM[926] = 23'h66ecd;
    RAM[927] = 23'h65d2a;
    RAM[928] = 23'h64b8a;
    RAM[929] = 23'h639f0;
    RAM[930] = 23'h6285a;
    RAM[931] = 23'h616c9;
    RAM[932] = 23'h6053c;
    RAM[933] = 23'h5f3b4;
    RAM[934] = 23'h5e231;
    RAM[935] = 23'h5d0b2;
    RAM[936] = 23'h5bf37;
    RAM[937] = 23'h5adc2;
    RAM[938] = 23'h59c50;
    RAM[939] = 23'h58ae4;
    RAM[940] = 23'h5797c;
    RAM[941] = 23'h56818;
    RAM[942] = 23'h556b9;
    RAM[943] = 23'h5455e;
    RAM[944] = 23'h53408;
    RAM[945] = 23'h522b7;
    RAM[946] = 23'h5116a;
    RAM[947] = 23'h50021;
    RAM[948] = 23'h4eedd;
    RAM[949] = 23'h4dd9e;
    RAM[950] = 23'h4cc63;
    RAM[951] = 23'h4bb2c;
    RAM[952] = 23'h4a9fa;
    RAM[953] = 23'h498cc;
    RAM[954] = 23'h487a3;
    RAM[955] = 23'h4767e;
    RAM[956] = 23'h4655e;
    RAM[957] = 23'h45442;
    RAM[958] = 23'h4432a;
    RAM[959] = 23'h43217;
    RAM[960] = 23'h42108;
    RAM[961] = 23'h40ffe;
    RAM[962] = 23'h3fef8;
    RAM[963] = 23'h3edf6;
    RAM[964] = 23'h3dcf9;
    RAM[965] = 23'h3cc00;
    RAM[966] = 23'h3bb0c;
    RAM[967] = 23'h3aa1c;
    RAM[968] = 23'h39930;
    RAM[969] = 23'h38849;
    RAM[970] = 23'h37766;
    RAM[971] = 23'h36687;
    RAM[972] = 23'h355ad;
    RAM[973] = 23'h344d7;
    RAM[974] = 23'h33405;
    RAM[975] = 23'h32338;
    RAM[976] = 23'h3126f;
    RAM[977] = 23'h301aa;
    RAM[978] = 23'h2f0e9;
    RAM[979] = 23'h2e02d;
    RAM[980] = 23'h2cf75;
    RAM[981] = 23'h2bec1;
    RAM[982] = 23'h2ae12;
    RAM[983] = 23'h29d67;
    RAM[984] = 23'h28cc0;
    RAM[985] = 23'h27c1d;
    RAM[986] = 23'h26b7f;
    RAM[987] = 23'h25ae4;
    RAM[988] = 23'h24a4e;
    RAM[989] = 23'h239bd;
    RAM[990] = 23'h2292f;
    RAM[991] = 23'h218a6;
    RAM[992] = 23'h20820;
    RAM[993] = 23'h1f7a0;
    RAM[994] = 23'h1e723;
    RAM[995] = 23'h1d6aa;
    RAM[996] = 23'h1c636;
    RAM[997] = 23'h1b5c5;
    RAM[998] = 23'h1a559;
    RAM[999] = 23'h194f1;
    RAM[1000] = 23'h1848e;
    RAM[1001] = 23'h1742e;
    RAM[1002] = 23'h163d2;
    RAM[1003] = 23'h1537b;
    RAM[1004] = 23'h14328;
    RAM[1005] = 23'h132d9;
    RAM[1006] = 23'h1228e;
    RAM[1007] = 23'h11247;
    RAM[1008] = 23'h10204;
    RAM[1009] = 23'hf1c5;
    RAM[1010] = 23'he18b;
    RAM[1011] = 23'hd154;
    RAM[1012] = 23'hc122;
    RAM[1013] = 23'hb0f3;
    RAM[1014] = 23'ha0c9;
    RAM[1015] = 23'h90a3;
    RAM[1016] = 23'h8080;
    RAM[1017] = 23'h7062;
    RAM[1018] = 23'h6048;
    RAM[1019] = 23'h5032;
    RAM[1020] = 23'h4020;
    RAM[1021] = 23'h3012;
    RAM[1022] = 23'h2008;
    RAM[1023] = 23'h1002;
    end
endmodule


module finv_grad_table (
    input wire clk, 
    input wire [9:0] addr,
    output reg [12:0] grd);

    reg [12:0] RAM [1023:0];
    always @(posedge clk)
        grd <= RAM[addr];
    initial begin
        RAM[0] = 13'h1ff8;
        RAM[1] = 13'h1fe8;
        RAM[2] = 13'h1fd8;
        RAM[3] = 13'h1fc8;
        RAM[4] = 13'h1fb8;
        RAM[5] = 13'h1fa8;
        RAM[6] = 13'h1f98;
        RAM[7] = 13'h1f89;
        RAM[8] = 13'h1f79;
        RAM[9] = 13'h1f6a;
        RAM[10] = 13'h1f5a;
        RAM[11] = 13'h1f4b;
        RAM[12] = 13'h1f3b;
        RAM[13] = 13'h1f2c;
        RAM[14] = 13'h1f1c;
        RAM[15] = 13'h1f0d;
        RAM[16] = 13'h1efe;
        RAM[17] = 13'h1eef;
        RAM[18] = 13'h1edf;
        RAM[19] = 13'h1ed0;
        RAM[20] = 13'h1ec1;
        RAM[21] = 13'h1eb2;
        RAM[22] = 13'h1ea3;
        RAM[23] = 13'h1e94;
        RAM[24] = 13'h1e85;
        RAM[25] = 13'h1e76;
        RAM[26] = 13'h1e67;
        RAM[27] = 13'h1e59;
        RAM[28] = 13'h1e4a;
        RAM[29] = 13'h1e3b;
        RAM[30] = 13'h1e2c;
        RAM[31] = 13'h1e1e;
        RAM[32] = 13'h1e0f;
        RAM[33] = 13'h1e01;
        RAM[34] = 13'h1df2;
        RAM[35] = 13'h1de4;
        RAM[36] = 13'h1dd5;
        RAM[37] = 13'h1dc7;
        RAM[38] = 13'h1db9;
        RAM[39] = 13'h1daa;
        RAM[40] = 13'h1d9c;
        RAM[41] = 13'h1d8e;
        RAM[42] = 13'h1d80;
        RAM[43] = 13'h1d71;
        RAM[44] = 13'h1d63;
        RAM[45] = 13'h1d55;
        RAM[46] = 13'h1d47;
        RAM[47] = 13'h1d39;
        RAM[48] = 13'h1d2b;
        RAM[49] = 13'h1d1d;
        RAM[50] = 13'h1d10;
        RAM[51] = 13'h1d02;
        RAM[52] = 13'h1cf4;
        RAM[53] = 13'h1ce6;
        RAM[54] = 13'h1cd8;
        RAM[55] = 13'h1ccb;
        RAM[56] = 13'h1cbd;
        RAM[57] = 13'h1cb0;
        RAM[58] = 13'h1ca2;
        RAM[59] = 13'h1c94;
        RAM[60] = 13'h1c87;
        RAM[61] = 13'h1c7a;
        RAM[62] = 13'h1c6c;
        RAM[63] = 13'h1c5f;
        RAM[64] = 13'h1c51;
        RAM[65] = 13'h1c44;
        RAM[66] = 13'h1c37;
        RAM[67] = 13'h1c2a;
        RAM[68] = 13'h1c1c;
        RAM[69] = 13'h1c0f;
        RAM[70] = 13'h1c02;
        RAM[71] = 13'h1bf5;
        RAM[72] = 13'h1be8;
        RAM[73] = 13'h1bdb;
        RAM[74] = 13'h1bce;
        RAM[75] = 13'h1bc1;
        RAM[76] = 13'h1bb4;
        RAM[77] = 13'h1ba7;
        RAM[78] = 13'h1b9a;
        RAM[79] = 13'h1b8e;
        RAM[80] = 13'h1b81;
        RAM[81] = 13'h1b74;
        RAM[82] = 13'h1b67;
        RAM[83] = 13'h1b5b;
        RAM[84] = 13'h1b4e;
        RAM[85] = 13'h1b42;
        RAM[86] = 13'h1b35;
        RAM[87] = 13'h1b28;
        RAM[88] = 13'h1b1c;
        RAM[89] = 13'h1b10;
        RAM[90] = 13'h1b03;
        RAM[91] = 13'h1af7;
        RAM[92] = 13'h1aea;
        RAM[93] = 13'h1ade;
        RAM[94] = 13'h1ad2;
        RAM[95] = 13'h1ac5;
        RAM[96] = 13'h1ab9;
        RAM[97] = 13'h1aad;
        RAM[98] = 13'h1aa1;
        RAM[99] = 13'h1a95;
        RAM[100] = 13'h1a89;
        RAM[101] = 13'h1a7d;
        RAM[102] = 13'h1a71;
        RAM[103] = 13'h1a65;
        RAM[104] = 13'h1a59;
        RAM[105] = 13'h1a4d;
        RAM[106] = 13'h1a41;
        RAM[107] = 13'h1a35;
        RAM[108] = 13'h1a29;
        RAM[109] = 13'h1a1d;
        RAM[110] = 13'h1a11;
        RAM[111] = 13'h1a06;
        RAM[112] = 13'h19fa;
        RAM[113] = 13'h19ee;
        RAM[114] = 13'h19e3;
        RAM[115] = 13'h19d7;
        RAM[116] = 13'h19cb;
        RAM[117] = 13'h19c0;
        RAM[118] = 13'h19b4;
        RAM[119] = 13'h19a9;
        RAM[120] = 13'h199d;
        RAM[121] = 13'h1992;
        RAM[122] = 13'h1986;
        RAM[123] = 13'h197b;
        RAM[124] = 13'h1970;
        RAM[125] = 13'h1964;
        RAM[126] = 13'h1959;
        RAM[127] = 13'h194e;
        RAM[128] = 13'h1943;
        RAM[129] = 13'h1937;
        RAM[130] = 13'h192c;
        RAM[131] = 13'h1921;
        RAM[132] = 13'h1916;
        RAM[133] = 13'h190b;
        RAM[134] = 13'h1900;
        RAM[135] = 13'h18f5;
        RAM[136] = 13'h18ea;
        RAM[137] = 13'h18df;
        RAM[138] = 13'h18d4;
        RAM[139] = 13'h18c9;
        RAM[140] = 13'h18be;
        RAM[141] = 13'h18b3;
        RAM[142] = 13'h18a8;
        RAM[143] = 13'h189d;
        RAM[144] = 13'h1893;
        RAM[145] = 13'h1888;
        RAM[146] = 13'h187d;
        RAM[147] = 13'h1873;
        RAM[148] = 13'h1868;
        RAM[149] = 13'h185d;
        RAM[150] = 13'h1853;
        RAM[151] = 13'h1848;
        RAM[152] = 13'h183d;
        RAM[153] = 13'h1833;
        RAM[154] = 13'h1828;
        RAM[155] = 13'h181e;
        RAM[156] = 13'h1813;
        RAM[157] = 13'h1809;
        RAM[158] = 13'h17ff;
        RAM[159] = 13'h17f4;
        RAM[160] = 13'h17ea;
        RAM[161] = 13'h17e0;
        RAM[162] = 13'h17d5;
        RAM[163] = 13'h17cb;
        RAM[164] = 13'h17c1;
        RAM[165] = 13'h17b7;
        RAM[166] = 13'h17ac;
        RAM[167] = 13'h17a2;
        RAM[168] = 13'h1798;
        RAM[169] = 13'h178e;
        RAM[170] = 13'h1784;
        RAM[171] = 13'h177a;
        RAM[172] = 13'h1770;
        RAM[173] = 13'h1766;
        RAM[174] = 13'h175c;
        RAM[175] = 13'h1752;
        RAM[176] = 13'h1748;
        RAM[177] = 13'h173e;
        RAM[178] = 13'h1734;
        RAM[179] = 13'h172a;
        RAM[180] = 13'h1720;
        RAM[181] = 13'h1716;
        RAM[182] = 13'h170d;
        RAM[183] = 13'h1703;
        RAM[184] = 13'h16f9;
        RAM[185] = 13'h16ef;
        RAM[186] = 13'h16e6;
        RAM[187] = 13'h16dc;
        RAM[188] = 13'h16d2;
        RAM[189] = 13'h16c9;
        RAM[190] = 13'h16bf;
        RAM[191] = 13'h16b6;
        RAM[192] = 13'h16ac;
        RAM[193] = 13'h16a2;
        RAM[194] = 13'h1699;
        RAM[195] = 13'h168f;
        RAM[196] = 13'h1686;
        RAM[197] = 13'h167d;
        RAM[198] = 13'h1673;
        RAM[199] = 13'h166a;
        RAM[200] = 13'h1660;
        RAM[201] = 13'h1657;
        RAM[202] = 13'h164e;
        RAM[203] = 13'h1644;
        RAM[204] = 13'h163b;
        RAM[205] = 13'h1632;
        RAM[206] = 13'h1629;
        RAM[207] = 13'h161f;
        RAM[208] = 13'h1616;
        RAM[209] = 13'h160d;
        RAM[210] = 13'h1604;
        RAM[211] = 13'h15fb;
        RAM[212] = 13'h15f2;
        RAM[213] = 13'h15e9;
        RAM[214] = 13'h15e0;
        RAM[215] = 13'h15d7;
        RAM[216] = 13'h15ce;
        RAM[217] = 13'h15c5;
        RAM[218] = 13'h15bc;
        RAM[219] = 13'h15b3;
        RAM[220] = 13'h15aa;
        RAM[221] = 13'h15a1;
        RAM[222] = 13'h1598;
        RAM[223] = 13'h158f;
        RAM[224] = 13'h1586;
        RAM[225] = 13'h157d;
        RAM[226] = 13'h1575;
        RAM[227] = 13'h156c;
        RAM[228] = 13'h1563;
        RAM[229] = 13'h155a;
        RAM[230] = 13'h1552;
        RAM[231] = 13'h1549;
        RAM[232] = 13'h1540;
        RAM[233] = 13'h1538;
        RAM[234] = 13'h152f;
        RAM[235] = 13'h1526;
        RAM[236] = 13'h151e;
        RAM[237] = 13'h1515;
        RAM[238] = 13'h150d;
        RAM[239] = 13'h1504;
        RAM[240] = 13'h14fc;
        RAM[241] = 13'h14f3;
        RAM[242] = 13'h14eb;
        RAM[243] = 13'h14e2;
        RAM[244] = 13'h14da;
        RAM[245] = 13'h14d1;
        RAM[246] = 13'h14c9;
        RAM[247] = 13'h14c1;
        RAM[248] = 13'h14b8;
        RAM[249] = 13'h14b0;
        RAM[250] = 13'h14a8;
        RAM[251] = 13'h149f;
        RAM[252] = 13'h1497;
        RAM[253] = 13'h148f;
        RAM[254] = 13'h1487;
        RAM[255] = 13'h147e;
        RAM[256] = 13'h1476;
        RAM[257] = 13'h146e;
        RAM[258] = 13'h1466;
        RAM[259] = 13'h145e;
        RAM[260] = 13'h1456;
        RAM[261] = 13'h144e;
        RAM[262] = 13'h1446;
        RAM[263] = 13'h143d;
        RAM[264] = 13'h1435;
        RAM[265] = 13'h142d;
        RAM[266] = 13'h1425;
        RAM[267] = 13'h141d;
        RAM[268] = 13'h1415;
        RAM[269] = 13'h140e;
        RAM[270] = 13'h1406;
        RAM[271] = 13'h13fe;
        RAM[272] = 13'h13f6;
        RAM[273] = 13'h13ee;
        RAM[274] = 13'h13e6;
        RAM[275] = 13'h13de;
        RAM[276] = 13'h13d6;
        RAM[277] = 13'h13cf;
        RAM[278] = 13'h13c7;
        RAM[279] = 13'h13bf;
        RAM[280] = 13'h13b7;
        RAM[281] = 13'h13b0;
        RAM[282] = 13'h13a8;
        RAM[283] = 13'h13a0;
        RAM[284] = 13'h1398;
        RAM[285] = 13'h1391;
        RAM[286] = 13'h1389;
        RAM[287] = 13'h1382;
        RAM[288] = 13'h137a;
        RAM[289] = 13'h1372;
        RAM[290] = 13'h136b;
        RAM[291] = 13'h1363;
        RAM[292] = 13'h135c;
        RAM[293] = 13'h1354;
        RAM[294] = 13'h134d;
        RAM[295] = 13'h1345;
        RAM[296] = 13'h133e;
        RAM[297] = 13'h1336;
        RAM[298] = 13'h132f;
        RAM[299] = 13'h1327;
        RAM[300] = 13'h1320;
        RAM[301] = 13'h1319;
        RAM[302] = 13'h1311;
        RAM[303] = 13'h130a;
        RAM[304] = 13'h1303;
        RAM[305] = 13'h12fb;
        RAM[306] = 13'h12f4;
        RAM[307] = 13'h12ed;
        RAM[308] = 13'h12e5;
        RAM[309] = 13'h12de;
        RAM[310] = 13'h12d7;
        RAM[311] = 13'h12d0;
        RAM[312] = 13'h12c8;
        RAM[313] = 13'h12c1;
        RAM[314] = 13'h12ba;
        RAM[315] = 13'h12b3;
        RAM[316] = 13'h12ac;
        RAM[317] = 13'h12a5;
        RAM[318] = 13'h129e;
        RAM[319] = 13'h1296;
        RAM[320] = 13'h128f;
        RAM[321] = 13'h1288;
        RAM[322] = 13'h1281;
        RAM[323] = 13'h127a;
        RAM[324] = 13'h1273;
        RAM[325] = 13'h126c;
        RAM[326] = 13'h1265;
        RAM[327] = 13'h125e;
        RAM[328] = 13'h1257;
        RAM[329] = 13'h1250;
        RAM[330] = 13'h124a;
        RAM[331] = 13'h1243;
        RAM[332] = 13'h123c;
        RAM[333] = 13'h1235;
        RAM[334] = 13'h122e;
        RAM[335] = 13'h1227;
        RAM[336] = 13'h1220;
        RAM[337] = 13'h1219;
        RAM[338] = 13'h1213;
        RAM[339] = 13'h120c;
        RAM[340] = 13'h1205;
        RAM[341] = 13'h11fe;
        RAM[342] = 13'h11f8;
        RAM[343] = 13'h11f1;
        RAM[344] = 13'h11ea;
        RAM[345] = 13'h11e4;
        RAM[346] = 13'h11dd;
        RAM[347] = 13'h11d6;
        RAM[348] = 13'h11d0;
        RAM[349] = 13'h11c9;
        RAM[350] = 13'h11c2;
        RAM[351] = 13'h11bc;
        RAM[352] = 13'h11b5;
        RAM[353] = 13'h11ae;
        RAM[354] = 13'h11a8;
        RAM[355] = 13'h11a1;
        RAM[356] = 13'h119b;
        RAM[357] = 13'h1194;
        RAM[358] = 13'h118e;
        RAM[359] = 13'h1187;
        RAM[360] = 13'h1181;
        RAM[361] = 13'h117a;
        RAM[362] = 13'h1174;
        RAM[363] = 13'h116d;
        RAM[364] = 13'h1167;
        RAM[365] = 13'h1161;
        RAM[366] = 13'h115a;
        RAM[367] = 13'h1154;
        RAM[368] = 13'h114d;
        RAM[369] = 13'h1147;
        RAM[370] = 13'h1141;
        RAM[371] = 13'h113a;
        RAM[372] = 13'h1134;
        RAM[373] = 13'h112e;
        RAM[374] = 13'h1128;
        RAM[375] = 13'h1121;
        RAM[376] = 13'h111b;
        RAM[377] = 13'h1115;
        RAM[378] = 13'h110f;
        RAM[379] = 13'h1108;
        RAM[380] = 13'h1102;
        RAM[381] = 13'h10fc;
        RAM[382] = 13'h10f6;
        RAM[383] = 13'h10f0;
        RAM[384] = 13'h10e9;
        RAM[385] = 13'h10e3;
        RAM[386] = 13'h10dd;
        RAM[387] = 13'h10d7;
        RAM[388] = 13'h10d1;
        RAM[389] = 13'h10cb;
        RAM[390] = 13'h10c5;
        RAM[391] = 13'h10bf;
        RAM[392] = 13'h10b9;
        RAM[393] = 13'h10b3;
        RAM[394] = 13'h10ad;
        RAM[395] = 13'h10a7;
        RAM[396] = 13'h10a1;
        RAM[397] = 13'h109b;
        RAM[398] = 13'h1095;
        RAM[399] = 13'h108f;
        RAM[400] = 13'h1089;
        RAM[401] = 13'h1083;
        RAM[402] = 13'h107d;
        RAM[403] = 13'h1077;
        RAM[404] = 13'h1071;
        RAM[405] = 13'h106b;
        RAM[406] = 13'h1065;
        RAM[407] = 13'h105f;
        RAM[408] = 13'h105a;
        RAM[409] = 13'h1054;
        RAM[410] = 13'h104e;
        RAM[411] = 13'h1048;
        RAM[412] = 13'h1042;
        RAM[413] = 13'h103c;
        RAM[414] = 13'h1037;
        RAM[415] = 13'h1031;
        RAM[416] = 13'h102b;
        RAM[417] = 13'h1025;
        RAM[418] = 13'h1020;
        RAM[419] = 13'h101a;
        RAM[420] = 13'h1014;
        RAM[421] = 13'h100f;
        RAM[422] = 13'h1009;
        RAM[423] = 13'h1003;
        RAM[424] = 13'hffe;
        RAM[425] = 13'hff8;
        RAM[426] = 13'hff2;
        RAM[427] = 13'hfed;
        RAM[428] = 13'hfe7;
        RAM[429] = 13'hfe1;
        RAM[430] = 13'hfdc;
        RAM[431] = 13'hfd6;
        RAM[432] = 13'hfd1;
        RAM[433] = 13'hfcb;
        RAM[434] = 13'hfc6;
        RAM[435] = 13'hfc0;
        RAM[436] = 13'hfbb;
        RAM[437] = 13'hfb5;
        RAM[438] = 13'hfb0;
        RAM[439] = 13'hfaa;
        RAM[440] = 13'hfa5;
        RAM[441] = 13'hf9f;
        RAM[442] = 13'hf9a;
        RAM[443] = 13'hf94;
        RAM[444] = 13'hf8f;
        RAM[445] = 13'hf89;
        RAM[446] = 13'hf84;
        RAM[447] = 13'hf7f;
        RAM[448] = 13'hf79;
        RAM[449] = 13'hf74;
        RAM[450] = 13'hf6e;
        RAM[451] = 13'hf69;
        RAM[452] = 13'hf64;
        RAM[453] = 13'hf5e;
        RAM[454] = 13'hf59;
        RAM[455] = 13'hf54;
        RAM[456] = 13'hf4e;
        RAM[457] = 13'hf49;
        RAM[458] = 13'hf44;
        RAM[459] = 13'hf3f;
        RAM[460] = 13'hf39;
        RAM[461] = 13'hf34;
        RAM[462] = 13'hf2f;
        RAM[463] = 13'hf2a;
        RAM[464] = 13'hf24;
        RAM[465] = 13'hf1f;
        RAM[466] = 13'hf1a;
        RAM[467] = 13'hf15;
        RAM[468] = 13'hf10;
        RAM[469] = 13'hf0b;
        RAM[470] = 13'hf05;
        RAM[471] = 13'hf00;
        RAM[472] = 13'hefb;
        RAM[473] = 13'hef6;
        RAM[474] = 13'hef1;
        RAM[475] = 13'heec;
        RAM[476] = 13'hee7;
        RAM[477] = 13'hee2;
        RAM[478] = 13'hedd;
        RAM[479] = 13'hed7;
        RAM[480] = 13'hed2;
        RAM[481] = 13'hecd;
        RAM[482] = 13'hec8;
        RAM[483] = 13'hec3;
        RAM[484] = 13'hebe;
        RAM[485] = 13'heb9;
        RAM[486] = 13'heb4;
        RAM[487] = 13'heaf;
        RAM[488] = 13'heaa;
        RAM[489] = 13'hea5;
        RAM[490] = 13'hea0;
        RAM[491] = 13'he9c;
        RAM[492] = 13'he97;
        RAM[493] = 13'he92;
        RAM[494] = 13'he8d;
        RAM[495] = 13'he88;
        RAM[496] = 13'he83;
        RAM[497] = 13'he7e;
        RAM[498] = 13'he79;
        RAM[499] = 13'he74;
        RAM[500] = 13'he70;
        RAM[501] = 13'he6b;
        RAM[502] = 13'he66;
        RAM[503] = 13'he61;
        RAM[504] = 13'he5c;
        RAM[505] = 13'he57;
        RAM[506] = 13'he53;
        RAM[507] = 13'he4e;
        RAM[508] = 13'he49;
        RAM[509] = 13'he44;
        RAM[510] = 13'he40;
        RAM[511] = 13'he3b;
        RAM[512] = 13'he36;
        RAM[513] = 13'he31;
        RAM[514] = 13'he2d;
        RAM[515] = 13'he28;
        RAM[516] = 13'he23;
        RAM[517] = 13'he1e;
        RAM[518] = 13'he1a;
        RAM[519] = 13'he15;
        RAM[520] = 13'he10;
        RAM[521] = 13'he0c;
        RAM[522] = 13'he07;
        RAM[523] = 13'he02;
        RAM[524] = 13'hdfe;
        RAM[525] = 13'hdf9;
        RAM[526] = 13'hdf5;
        RAM[527] = 13'hdf0;
        RAM[528] = 13'hdeb;
        RAM[529] = 13'hde7;
        RAM[530] = 13'hde2;
        RAM[531] = 13'hdde;
        RAM[532] = 13'hdd9;
        RAM[533] = 13'hdd5;
        RAM[534] = 13'hdd0;
        RAM[535] = 13'hdcb;
        RAM[536] = 13'hdc7;
        RAM[537] = 13'hdc2;
        RAM[538] = 13'hdbe;
        RAM[539] = 13'hdb9;
        RAM[540] = 13'hdb5;
        RAM[541] = 13'hdb0;
        RAM[542] = 13'hdac;
        RAM[543] = 13'hda8;
        RAM[544] = 13'hda3;
        RAM[545] = 13'hd9f;
        RAM[546] = 13'hd9a;
        RAM[547] = 13'hd96;
        RAM[548] = 13'hd91;
        RAM[549] = 13'hd8d;
        RAM[550] = 13'hd89;
        RAM[551] = 13'hd84;
        RAM[552] = 13'hd80;
        RAM[553] = 13'hd7b;
        RAM[554] = 13'hd77;
        RAM[555] = 13'hd73;
        RAM[556] = 13'hd6e;
        RAM[557] = 13'hd6a;
        RAM[558] = 13'hd66;
        RAM[559] = 13'hd61;
        RAM[560] = 13'hd5d;
        RAM[561] = 13'hd59;
        RAM[562] = 13'hd54;
        RAM[563] = 13'hd50;
        RAM[564] = 13'hd4c;
        RAM[565] = 13'hd47;
        RAM[566] = 13'hd43;
        RAM[567] = 13'hd3f;
        RAM[568] = 13'hd3b;
        RAM[569] = 13'hd36;
        RAM[570] = 13'hd32;
        RAM[571] = 13'hd2e;
        RAM[572] = 13'hd2a;
        RAM[573] = 13'hd25;
        RAM[574] = 13'hd21;
        RAM[575] = 13'hd1d;
        RAM[576] = 13'hd19;
        RAM[577] = 13'hd15;
        RAM[578] = 13'hd10;
        RAM[579] = 13'hd0c;
        RAM[580] = 13'hd08;
        RAM[581] = 13'hd04;
        RAM[582] = 13'hd00;
        RAM[583] = 13'hcfc;
        RAM[584] = 13'hcf8;
        RAM[585] = 13'hcf3;
        RAM[586] = 13'hcef;
        RAM[587] = 13'hceb;
        RAM[588] = 13'hce7;
        RAM[589] = 13'hce3;
        RAM[590] = 13'hcdf;
        RAM[591] = 13'hcdb;
        RAM[592] = 13'hcd7;
        RAM[593] = 13'hcd3;
        RAM[594] = 13'hccf;
        RAM[595] = 13'hccb;
        RAM[596] = 13'hcc7;
        RAM[597] = 13'hcc3;
        RAM[598] = 13'hcbf;
        RAM[599] = 13'hcbb;
        RAM[600] = 13'hcb6;
        RAM[601] = 13'hcb2;
        RAM[602] = 13'hcae;
        RAM[603] = 13'hcab;
        RAM[604] = 13'hca7;
        RAM[605] = 13'hca3;
        RAM[606] = 13'hc9f;
        RAM[607] = 13'hc9b;
        RAM[608] = 13'hc97;
        RAM[609] = 13'hc93;
        RAM[610] = 13'hc8f;
        RAM[611] = 13'hc8b;
        RAM[612] = 13'hc87;
        RAM[613] = 13'hc83;
        RAM[614] = 13'hc7f;
        RAM[615] = 13'hc7b;
        RAM[616] = 13'hc77;
        RAM[617] = 13'hc73;
        RAM[618] = 13'hc70;
        RAM[619] = 13'hc6c;
        RAM[620] = 13'hc68;
        RAM[621] = 13'hc64;
        RAM[622] = 13'hc60;
        RAM[623] = 13'hc5c;
        RAM[624] = 13'hc58;
        RAM[625] = 13'hc55;
        RAM[626] = 13'hc51;
        RAM[627] = 13'hc4d;
        RAM[628] = 13'hc49;
        RAM[629] = 13'hc45;
        RAM[630] = 13'hc42;
        RAM[631] = 13'hc3e;
        RAM[632] = 13'hc3a;
        RAM[633] = 13'hc36;
        RAM[634] = 13'hc32;
        RAM[635] = 13'hc2f;
        RAM[636] = 13'hc2b;
        RAM[637] = 13'hc27;
        RAM[638] = 13'hc23;
        RAM[639] = 13'hc20;
        RAM[640] = 13'hc1c;
        RAM[641] = 13'hc18;
        RAM[642] = 13'hc14;
        RAM[643] = 13'hc11;
        RAM[644] = 13'hc0d;
        RAM[645] = 13'hc09;
        RAM[646] = 13'hc06;
        RAM[647] = 13'hc02;
        RAM[648] = 13'hbfe;
        RAM[649] = 13'hbfb;
        RAM[650] = 13'hbf7;
        RAM[651] = 13'hbf3;
        RAM[652] = 13'hbf0;
        RAM[653] = 13'hbec;
        RAM[654] = 13'hbe8;
        RAM[655] = 13'hbe5;
        RAM[656] = 13'hbe1;
        RAM[657] = 13'hbde;
        RAM[658] = 13'hbda;
        RAM[659] = 13'hbd6;
        RAM[660] = 13'hbd3;
        RAM[661] = 13'hbcf;
        RAM[662] = 13'hbcc;
        RAM[663] = 13'hbc8;
        RAM[664] = 13'hbc4;
        RAM[665] = 13'hbc1;
        RAM[666] = 13'hbbd;
        RAM[667] = 13'hbba;
        RAM[668] = 13'hbb6;
        RAM[669] = 13'hbb3;
        RAM[670] = 13'hbaf;
        RAM[671] = 13'hbac;
        RAM[672] = 13'hba8;
        RAM[673] = 13'hba5;
        RAM[674] = 13'hba1;
        RAM[675] = 13'hb9e;
        RAM[676] = 13'hb9a;
        RAM[677] = 13'hb97;
        RAM[678] = 13'hb93;
        RAM[679] = 13'hb90;
        RAM[680] = 13'hb8c;
        RAM[681] = 13'hb89;
        RAM[682] = 13'hb85;
        RAM[683] = 13'hb82;
        RAM[684] = 13'hb7e;
        RAM[685] = 13'hb7b;
        RAM[686] = 13'hb77;
        RAM[687] = 13'hb74;
        RAM[688] = 13'hb71;
        RAM[689] = 13'hb6d;
        RAM[690] = 13'hb6a;
        RAM[691] = 13'hb66;
        RAM[692] = 13'hb63;
        RAM[693] = 13'hb60;
        RAM[694] = 13'hb5c;
        RAM[695] = 13'hb59;
        RAM[696] = 13'hb55;
        RAM[697] = 13'hb52;
        RAM[698] = 13'hb4f;
        RAM[699] = 13'hb4b;
        RAM[700] = 13'hb48;
        RAM[701] = 13'hb45;
        RAM[702] = 13'hb41;
        RAM[703] = 13'hb3e;
        RAM[704] = 13'hb3b;
        RAM[705] = 13'hb37;
        RAM[706] = 13'hb34;
        RAM[707] = 13'hb31;
        RAM[708] = 13'hb2d;
        RAM[709] = 13'hb2a;
        RAM[710] = 13'hb27;
        RAM[711] = 13'hb23;
        RAM[712] = 13'hb20;
        RAM[713] = 13'hb1d;
        RAM[714] = 13'hb1a;
        RAM[715] = 13'hb16;
        RAM[716] = 13'hb13;
        RAM[717] = 13'hb10;
        RAM[718] = 13'hb0d;
        RAM[719] = 13'hb09;
        RAM[720] = 13'hb06;
        RAM[721] = 13'hb03;
        RAM[722] = 13'hb00;
        RAM[723] = 13'hafc;
        RAM[724] = 13'haf9;
        RAM[725] = 13'haf6;
        RAM[726] = 13'haf3;
        RAM[727] = 13'haf0;
        RAM[728] = 13'haec;
        RAM[729] = 13'hae9;
        RAM[730] = 13'hae6;
        RAM[731] = 13'hae3;
        RAM[732] = 13'hae0;
        RAM[733] = 13'hadc;
        RAM[734] = 13'had9;
        RAM[735] = 13'had6;
        RAM[736] = 13'had3;
        RAM[737] = 13'had0;
        RAM[738] = 13'hacd;
        RAM[739] = 13'haca;
        RAM[740] = 13'hac6;
        RAM[741] = 13'hac3;
        RAM[742] = 13'hac0;
        RAM[743] = 13'habd;
        RAM[744] = 13'haba;
        RAM[745] = 13'hab7;
        RAM[746] = 13'hab4;
        RAM[747] = 13'hab1;
        RAM[748] = 13'haae;
        RAM[749] = 13'haab;
        RAM[750] = 13'haa7;
        RAM[751] = 13'haa4;
        RAM[752] = 13'haa1;
        RAM[753] = 13'ha9e;
        RAM[754] = 13'ha9b;
        RAM[755] = 13'ha98;
        RAM[756] = 13'ha95;
        RAM[757] = 13'ha92;
        RAM[758] = 13'ha8f;
        RAM[759] = 13'ha8c;
        RAM[760] = 13'ha89;
        RAM[761] = 13'ha86;
        RAM[762] = 13'ha83;
        RAM[763] = 13'ha80;
        RAM[764] = 13'ha7d;
        RAM[765] = 13'ha7a;
        RAM[766] = 13'ha77;
        RAM[767] = 13'ha74;
        RAM[768] = 13'ha71;
        RAM[769] = 13'ha6e;
        RAM[770] = 13'ha6b;
        RAM[771] = 13'ha68;
        RAM[772] = 13'ha65;
        RAM[773] = 13'ha62;
        RAM[774] = 13'ha5f;
        RAM[775] = 13'ha5c;
        RAM[776] = 13'ha59;
        RAM[777] = 13'ha56;
        RAM[778] = 13'ha53;
        RAM[779] = 13'ha50;
        RAM[780] = 13'ha4e;
        RAM[781] = 13'ha4b;
        RAM[782] = 13'ha48;
        RAM[783] = 13'ha45;
        RAM[784] = 13'ha42;
        RAM[785] = 13'ha3f;
        RAM[786] = 13'ha3c;
        RAM[787] = 13'ha39;
        RAM[788] = 13'ha36;
        RAM[789] = 13'ha33;
        RAM[790] = 13'ha31;
        RAM[791] = 13'ha2e;
        RAM[792] = 13'ha2b;
        RAM[793] = 13'ha28;
        RAM[794] = 13'ha25;
        RAM[795] = 13'ha22;
        RAM[796] = 13'ha1f;
        RAM[797] = 13'ha1c;
        RAM[798] = 13'ha1a;
        RAM[799] = 13'ha17;
        RAM[800] = 13'ha14;
        RAM[801] = 13'ha11;
        RAM[802] = 13'ha0e;
        RAM[803] = 13'ha0c;
        RAM[804] = 13'ha09;
        RAM[805] = 13'ha06;
        RAM[806] = 13'ha03;
        RAM[807] = 13'ha00;
        RAM[808] = 13'h9fe;
        RAM[809] = 13'h9fb;
        RAM[810] = 13'h9f8;
        RAM[811] = 13'h9f5;
        RAM[812] = 13'h9f2;
        RAM[813] = 13'h9f0;
        RAM[814] = 13'h9ed;
        RAM[815] = 13'h9ea;
        RAM[816] = 13'h9e7;
        RAM[817] = 13'h9e5;
        RAM[818] = 13'h9e2;
        RAM[819] = 13'h9df;
        RAM[820] = 13'h9dc;
        RAM[821] = 13'h9da;
        RAM[822] = 13'h9d7;
        RAM[823] = 13'h9d4;
        RAM[824] = 13'h9d1;
        RAM[825] = 13'h9cf;
        RAM[826] = 13'h9cc;
        RAM[827] = 13'h9c9;
        RAM[828] = 13'h9c7;
        RAM[829] = 13'h9c4;
        RAM[830] = 13'h9c1;
        RAM[831] = 13'h9be;
        RAM[832] = 13'h9bc;
        RAM[833] = 13'h9b9;
        RAM[834] = 13'h9b6;
        RAM[835] = 13'h9b4;
        RAM[836] = 13'h9b1;
        RAM[837] = 13'h9ae;
        RAM[838] = 13'h9ac;
        RAM[839] = 13'h9a9;
        RAM[840] = 13'h9a6;
        RAM[841] = 13'h9a4;
        RAM[842] = 13'h9a1;
        RAM[843] = 13'h99f;
        RAM[844] = 13'h99c;
        RAM[845] = 13'h999;
        RAM[846] = 13'h997;
        RAM[847] = 13'h994;
        RAM[848] = 13'h991;
        RAM[849] = 13'h98f;
        RAM[850] = 13'h98c;
        RAM[851] = 13'h98a;
        RAM[852] = 13'h987;
        RAM[853] = 13'h984;
        RAM[854] = 13'h982;
        RAM[855] = 13'h97f;
        RAM[856] = 13'h97d;
        RAM[857] = 13'h97a;
        RAM[858] = 13'h977;
        RAM[859] = 13'h975;
        RAM[860] = 13'h972;
        RAM[861] = 13'h970;
        RAM[862] = 13'h96d;
        RAM[863] = 13'h96b;
        RAM[864] = 13'h968;
        RAM[865] = 13'h966;
        RAM[866] = 13'h963;
        RAM[867] = 13'h960;
        RAM[868] = 13'h95e;
        RAM[869] = 13'h95b;
        RAM[870] = 13'h959;
        RAM[871] = 13'h956;
        RAM[872] = 13'h954;
        RAM[873] = 13'h951;
        RAM[874] = 13'h94f;
        RAM[875] = 13'h94c;
        RAM[876] = 13'h94a;
        RAM[877] = 13'h947;
        RAM[878] = 13'h945;
        RAM[879] = 13'h942;
        RAM[880] = 13'h940;
        RAM[881] = 13'h93d;
        RAM[882] = 13'h93b;
        RAM[883] = 13'h938;
        RAM[884] = 13'h936;
        RAM[885] = 13'h933;
        RAM[886] = 13'h931;
        RAM[887] = 13'h92e;
        RAM[888] = 13'h92c;
        RAM[889] = 13'h92a;
        RAM[890] = 13'h927;
        RAM[891] = 13'h925;
        RAM[892] = 13'h922;
        RAM[893] = 13'h920;
        RAM[894] = 13'h91d;
        RAM[895] = 13'h91b;
        RAM[896] = 13'h918;
        RAM[897] = 13'h916;
        RAM[898] = 13'h914;
        RAM[899] = 13'h911;
        RAM[900] = 13'h90f;
        RAM[901] = 13'h90c;
        RAM[902] = 13'h90a;
        RAM[903] = 13'h908;
        RAM[904] = 13'h905;
        RAM[905] = 13'h903;
        RAM[906] = 13'h900;
        RAM[907] = 13'h8fe;
        RAM[908] = 13'h8fc;
        RAM[909] = 13'h8f9;
        RAM[910] = 13'h8f7;
        RAM[911] = 13'h8f4;
        RAM[912] = 13'h8f2;
        RAM[913] = 13'h8f0;
        RAM[914] = 13'h8ed;
        RAM[915] = 13'h8eb;
        RAM[916] = 13'h8e9;
        RAM[917] = 13'h8e6;
        RAM[918] = 13'h8e4;
        RAM[919] = 13'h8e2;
        RAM[920] = 13'h8df;
        RAM[921] = 13'h8dd;
        RAM[922] = 13'h8db;
        RAM[923] = 13'h8d8;
        RAM[924] = 13'h8d6;
        RAM[925] = 13'h8d4;
        RAM[926] = 13'h8d1;
        RAM[927] = 13'h8cf;
        RAM[928] = 13'h8cd;
        RAM[929] = 13'h8ca;
        RAM[930] = 13'h8c8;
        RAM[931] = 13'h8c6;
        RAM[932] = 13'h8c4;
        RAM[933] = 13'h8c1;
        RAM[934] = 13'h8bf;
        RAM[935] = 13'h8bd;
        RAM[936] = 13'h8ba;
        RAM[937] = 13'h8b8;
        RAM[938] = 13'h8b6;
        RAM[939] = 13'h8b4;
        RAM[940] = 13'h8b1;
        RAM[941] = 13'h8af;
        RAM[942] = 13'h8ad;
        RAM[943] = 13'h8ab;
        RAM[944] = 13'h8a8;
        RAM[945] = 13'h8a6;
        RAM[946] = 13'h8a4;
        RAM[947] = 13'h8a2;
        RAM[948] = 13'h89f;
        RAM[949] = 13'h89d;
        RAM[950] = 13'h89b;
        RAM[951] = 13'h899;
        RAM[952] = 13'h896;
        RAM[953] = 13'h894;
        RAM[954] = 13'h892;
        RAM[955] = 13'h890;
        RAM[956] = 13'h88d;
        RAM[957] = 13'h88b;
        RAM[958] = 13'h889;
        RAM[959] = 13'h887;
        RAM[960] = 13'h885;
        RAM[961] = 13'h882;
        RAM[962] = 13'h880;
        RAM[963] = 13'h87e;
        RAM[964] = 13'h87c;
        RAM[965] = 13'h87a;
        RAM[966] = 13'h878;
        RAM[967] = 13'h875;
        RAM[968] = 13'h873;
        RAM[969] = 13'h871;
        RAM[970] = 13'h86f;
        RAM[971] = 13'h86d;
        RAM[972] = 13'h86b;
        RAM[973] = 13'h868;
        RAM[974] = 13'h866;
        RAM[975] = 13'h864;
        RAM[976] = 13'h862;
        RAM[977] = 13'h860;
        RAM[978] = 13'h85e;
        RAM[979] = 13'h85b;
        RAM[980] = 13'h859;
        RAM[981] = 13'h857;
        RAM[982] = 13'h855;
        RAM[983] = 13'h853;
        RAM[984] = 13'h851;
        RAM[985] = 13'h84f;
        RAM[986] = 13'h84d;
        RAM[987] = 13'h84a;
        RAM[988] = 13'h848;
        RAM[989] = 13'h846;
        RAM[990] = 13'h844;
        RAM[991] = 13'h842;
        RAM[992] = 13'h840;
        RAM[993] = 13'h83e;
        RAM[994] = 13'h83c;
        RAM[995] = 13'h83a;
        RAM[996] = 13'h838;
        RAM[997] = 13'h836;
        RAM[998] = 13'h833;
        RAM[999] = 13'h831;
        RAM[1000] = 13'h82f;
        RAM[1001] = 13'h82d;
        RAM[1002] = 13'h82b;
        RAM[1003] = 13'h829;
        RAM[1004] = 13'h827;
        RAM[1005] = 13'h825;
        RAM[1006] = 13'h823;
        RAM[1007] = 13'h821;
        RAM[1008] = 13'h81f;
        RAM[1009] = 13'h81d;
        RAM[1010] = 13'h81b;
        RAM[1011] = 13'h819;
        RAM[1012] = 13'h817;
        RAM[1013] = 13'h815;
        RAM[1014] = 13'h813;
        RAM[1015] = 13'h811;
        RAM[1016] = 13'h80f;
        RAM[1017] = 13'h80d;
        RAM[1018] = 13'h80b;
        RAM[1019] = 13'h809;
        RAM[1020] = 13'h807;
        RAM[1021] = 13'h805;
        RAM[1022] = 13'h803;
        RAM[1023] = 13'h801;
    end
 endmodule
`default_nettype wire
